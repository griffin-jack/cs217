
//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Thu Jan 15 14:27:17 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [168:0] this_dat;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [127:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_dat[127:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_dat[151:128];
  wire  nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_dat[168];
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd128)) data_data_rsci (
      .d(nl_data_data_rsci_d[127:0]),
      .z(data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d),
      .z(data_rw_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd153),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [168:0] this_dat;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Thu Jan 15 14:27:12 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [137:0] this_dat;
  output [127:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [127:0] nl_data_data_data_rsci_d;
  assign nl_data_data_data_rsci_d = this_dat[127:0];
  wire [7:0] nl_data_logical_addr_rsci_d;
  assign nl_data_logical_addr_rsci_d = this_dat[137:130];
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd7),
  .width(32'sd128)) data_data_data_rsci (
      .d(nl_data_data_data_rsci_d[127:0]),
      .z(data_data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd9),
  .width(32'sd8)) data_logical_addr_rsci (
      .d(nl_data_logical_addr_rsci_d[7:0]),
      .z(data_logical_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd11),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd152),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [137:0] this_dat;
  output [127:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_data_rsc_z(data_data_data_rsc_z),
      .data_logical_addr_rsc_z(data_logical_addr_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Wed Jan 14 11:37:19 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [255:0] this_dat;
  reg [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [255:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd13),
  .width(32'sd256)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd151),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd155)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Wed Jan 14 11:37:16 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd15),
  .width(32'sd1)) data_rsci (
      .d(this_dat),
      .z(data_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd17),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd150),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Thu Jan 15 14:27:15 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [127:0] this_dat;
  reg [127:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [127:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd18),
  .width(32'sd128)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd149),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd154)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [127:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module PECore_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // spyglass disable SYNTH_5121,W240
    input                s_rst;  // spyglass disable SYNTH_5121,W240
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a; //spyglass disable FlopEConst
                b_reg[0] <= b; //spyglass disable FlopEConst
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> ./PECore_mgc_muladd1_beh.v 
//muladd1
module PECore_mgc_muladd1(a,b,c,cst,d,z);
  // operation is z = a * (b + d) + c + cst
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_cst = 0;
  parameter signd_cst = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_axb = 1;
  parameter add_c = 1;
  parameter add_d = 1;
  parameter use_const = 1;

  function integer is_square_op;
    input integer alen;
  begin
    if (alen > 1) is_square_op = 0;
    else       is_square_op = 1;
  end endfunction

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_cst-1:0] cst; // spyglass disable SYNTH_5121,W240
  input  [width_d-1:0] d;
  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa;
  reg [width_b-signd_b:0] bb;
  reg [width_c-signd_c:0] cc;
  reg [width_d-signd_d:0] dd;
  reg [width_cst-signd_cst:0] cstin;

  localparam width_bd = (width_d) ? 1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b
                                                                          : width_d - signd_d)
                                  : width_b - signd_b;
  localparam is_square = is_square_op(width_a);
  localparam axb_len = (is_square)?width_bd+1+width_bd+1:width_a-signd_a+1+width_bd+1;

  reg [width_bd:0] bd;
  reg [axb_len-1:0] axb;



  // make all inputs signed
  always @(*) aa = signd_a ? a : {1'b0, a};
  always @(*) bb = signd_b ? b : {1'b0, b};
  generate if (width_c != 0) begin
    always @(*) cc = signd_c ? c : {1'b0, c};
  end endgenerate

  generate if (width_d) begin
    if ( !is_square) begin
      (* keep ="true" *) reg [width_d-signd_d:0] d_keep;
      always @(*) d_keep = signd_d ? d : {1'b0, d};
      always @(*) dd = d_keep;
    end else begin
      always @(*) dd = signd_d ? d : {1'b0, d};
    end
  end endgenerate

  always @(*) cstin = signd_cst ? cst : {1'b0, cst};

  // perform pre-adder
  generate
    if (width_d != 0) begin
      if (add_d) begin always @(*)  bd = $signed(bb) + $signed(dd); end
      else       begin always @(*)  bd = $signed(bb) - $signed(dd); end
    end else     begin always @(*)  bd = $signed(bb); end
  endgenerate

  generate
    if (is_square)
      always @(*) axb = $signed(bd) * $signed(bd);
    else
      always @(*) axb = $signed(aa) * $signed(bd);
  endgenerate

  // perform muladd1
  wire [width_z-1:0]  zz;

  generate
    if (use_const) begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc) + $signed(cstin); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc) + $signed(cstin); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb) + $signed(cstin); end else
      if (!add_axb && !add_c && width_c) begin assign zz = $signed(cstin) - $signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb) + $signed(cstin); end else
                                         begin assign zz = $signed(cstin) - $signed(axb); end
    end  else begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb); end else
      if (!add_axb && !add_c && width_c) begin assign zz = -$signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb); end else
                                         begin assign zz = -$signed(axb); end
    end
  endgenerate

  // adjust output
  assign z = zz;
endmodule // mgc_muladd1

//------> ./PECore_mgc_shift_l_beh_v5.v 
module PECore_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./PECore_mgc_mulacc_pipe_beh.v 
//mulacc
module PECore_mgc_mulacc_pipe(a,b,c,d,load,datavalid,clk,en,a_rst,s_rst,z);

  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_d = 1;
  parameter is_square = 0;
  parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
  parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
  parameter    a_rst_active =  1'b1;  // unused
  parameter    s_rst_active =  1'b1;  // unused
  parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
  parameter integer n_inreg = 32'd0;  // number of input registers

  function integer max_len;
    input integer a, b;
  begin
    if (a > b) max_len = a;
    else       max_len = b;
  end endfunction

  function integer min_len;
    input integer a, b;
  begin
    if (a > b) min_len = b;
    else       min_len = a;
  end endfunction

  localparam axb_stages = (stages>2) ? 1 : 0;

  localparam preadd_stages = (n_inreg>1) ? 1 : 0;
  localparam bb_stages = n_inreg - preadd_stages;
  localparam cc_stages = n_inreg + axb_stages;
  localparam cc_len = min_len(width_c-signd_c+1, width_z);

  localparam zz_stages = stages - axb_stages;

  localparam width_bd = (width_d>0) ? (1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b : width_d - signd_d)) : width_b - signd_b;
  localparam axb_len = (is_square)?width_bd+1+width_bd+1:width_a-signd_a+1+width_bd+1;

  localparam zz_len = max_len(axb_len, max_len(cc_len, width_z));

  reg [width_bd:0] bd [preadd_stages:0];

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_d-1:0] d; // spyglass disable SYNTH_5121,W240
  input                load;
  input                datavalid;

  input                clk;    // clock
  input                en;     // enable
  input                a_rst;  // spyglass disable SYNTH_5121,W240
  input                s_rst;  // spyglass disable SYNTH_5121,W240

  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa [n_inreg:0];
  reg [width_b-signd_b:0] bb [n_inreg:0];
  reg [width_c-signd_c:0] cc [cc_stages:0];
  reg [width_d-signd_d:0] dd [bb_stages:0];
  reg                     accum [cc_stages:0];
  reg                     vl [cc_stages:0];

  genvar i;

  // make all inputs signed
  always @(*) aa[n_inreg]   = signd_a ? a : {1'b0, a};
  always @(*) bb[bb_stages]   = signd_b ? b : {1'b0, b};
  generate if (width_d>0) begin
    always @(*) dd[bb_stages]   = signd_d ? d : {1'b0, d};
  end endgenerate
  always @(*) cc[cc_stages] = (signd_c | width_c >= width_z) ? c : {1'b0, c};
  always @(*) accum[cc_stages] = !load;
  always @(*) vl[cc_stages] = datavalid;

  // input registers
  generate if (n_inreg>0) begin
  for(i = n_inreg-1; i >= 0; i=i-1) begin:ab_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (bb_stages>0) begin
  for(i = bb_stages-1; i >= 0; i=i-1) begin:in_pipe_bd
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];
      if (width_d>0) begin  always @(posedge(clk)) if (en == enable_active) dd[i] <= dd[i+1]; end //spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];
      if (width_d>0) begin  always @(negedge(clk)) if (en == enable_active) dd[i] <= dd[i+1]; end //spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (cc_stages>0) begin
  for(i = cc_stages-1; i >= 0; i=i-1) begin:c_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) accum[i] <= accum[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) vl[i] <= vl[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) accum[i] <= accum[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) vl[i] <= vl[i+1];
    end
  end end endgenerate

  // perform pre-adder
  generate
    if (width_d>0) begin
      if (add_d != 0) begin always @(*)  bd[preadd_stages] = $signed(bb[0]) + $signed(dd[0]); end
      else            begin always @(*)  bd[preadd_stages] = $signed(bb[0]) - $signed(dd[0]); end
    end else          begin always @(*)  bd[preadd_stages] = $signed(bb[0]); end
  endgenerate
  generate if (preadd_stages>0) begin
  for(i = preadd_stages-1; i >= 0; i=i-1) begin:preadd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bd[i] <= bd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bd[i] <= bd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // perform muladd1
  reg [zz_len-1:0]  zz[zz_stages-1:0];
  wire [zz_len-1:0] z_or_c;
  reg [axb_len-1:0] axb[axb_stages:0];
  generate
    if (is_square>0)
      always @(*) axb[axb_stages] = $signed(bd[0]) * $signed(bd[0]);
    else
      always @(*) axb[axb_stages] = $signed(aa[0]) * $signed(bd[0]);
  endgenerate

  generate if (axb_stages>0) begin
  for(i = axb_stages-1; i >= 0; i=i-1) begin:axb_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  assign z_or_c = accum[0] ? $signed(zz[zz_stages-2]): $signed(cc[0]);
  always @(*) zz[zz_stages-1] = $signed(axb[0]) + $signed(z_or_c);

  // Output registers:
  generate for(i = zz_stages-2; i >= 0; i=i-1) begin:out_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active && (vl[0] || i != zz_stages-2)) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active && (vl[0] || i != zz_stages-2)) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end
  end endgenerate

  // adjust output
  // use a tmp var to satisfy W164a lint violations
  wire [width_z-1:0] z_out_tmp;
  assign z_out_tmp = zz[0][width_z-1:0];
  assign z = z_out_tmp;

endmodule // mgc_mulacc_pipe

//------> ./PECore_mgc_mul4acc_pipe_beh.v 
//mulacc
module PECore_mgc_mul4acc_pipe(a0,a1,b0,b1,c0,c1,d0,d1,e,load,datavalid,clk,en,a_rst,s_rst,z);

  parameter width_a0 = 0;
  parameter signd_a0 = 0;
  parameter width_a1 = 0;
  parameter signd_a1 = 0;
  parameter width_b0 = 0;
  parameter signd_b0 = 0;
  parameter width_b1 = 0;
  parameter signd_b1 = 0;
  parameter width_c0 = 0;
  parameter signd_c0 = 0;
  parameter width_c1 = 0;
  parameter signd_c1 = 0;
  parameter width_d0 = 0;
  parameter signd_d0 = 0;
  parameter width_d1 = 0;
  parameter signd_d1 = 0;
  parameter width_e  = 0;
  parameter signd_e  = 0;
  parameter width_z = 0;
  parameter add_a    = 1;
  parameter add_b    = 1;
  parameter add_c    = 1;
  parameter min_fb_size    = -1;

  parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
  parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
  parameter    a_rst_active =  1'b1;  // unused
  parameter    s_rst_active =  1'b1;  // unused
  parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
  parameter integer n_inreg = 32'd0;  // number of input registers

  function integer max_len;
    input integer a, b;
  begin
    if (a > b) max_len = a;
    else       max_len = b;
  end endfunction

  function integer min_len;
    input integer a, b;
  begin
    if (a > b) min_len = b;
    else       min_len = a;
  end endfunction

  localparam nb_prod_reg = 0;
  localparam nb_in_reg = n_inreg - nb_prod_reg;
  localparam nb_sop_reg = (stages>2)?1:0;
  localparam out_stages = stages - nb_sop_reg;

  localparam ee_len = min_len(width_e-signd_e+1, width_z);
  localparam zz_len = (min_fb_size>width_z)?min_fb_size:width_z;
  localparam proda_len = width_a0-signd_a0+width_a1-signd_a1+2;
  localparam prodb_len = width_b0-signd_b0+width_b1-signd_b1+2;
  localparam prodc_len = width_c0-signd_c0+width_c1-signd_c1+2;
  localparam prodd_len = width_d0-signd_d0+width_d1-signd_d1+2;
  localparam sop_len = 2 + max_len(proda_len,max_len(prodb_len,max_len(prodc_len,prodd_len)));

  localparam proda_pol  = (add_a>0)?1:-1;
  localparam prodb_pol  = (add_b>0)?1:-1;
  localparam prodc_pol  = (add_c>0)?1:-1;
  localparam prodd_pol  = 1;

  input  [width_a0-1:0] a0;
  input  [width_a1-1:0] a1;
  input  [width_b0-1:0] b0;
  input  [width_b1-1:0] b1;
  input  [width_c0-1:0] c0;
  input  [width_c1-1:0] c1;
  input  [width_d0-1:0] d0; // spyglass disable SYNTH_5121,W240
  input  [width_d1-1:0] d1; // spyglass disable SYNTH_5121,W240
  input  [width_e-1:0]  e;
  input                load;
  input                datavalid;

  input                clk;    // clock
  input                en;     // enable
  input                a_rst;  // spyglass disable SYNTH_5121,W240
  input                s_rst;  // spyglass disable SYNTH_5121,W240

  output [width_z-1:0] z;



  reg [width_a0-signd_a0:0] aa0 [nb_in_reg:0];
  reg [width_b0-signd_b0:0] bb0 [nb_in_reg:0];
  reg [width_c0-signd_c0:0] cc0 [nb_in_reg:0];
  reg [width_d0-signd_d0:0] dd0 [nb_in_reg:0];
  reg [width_a1-signd_a1:0] aa1 [nb_in_reg:0];
  reg [width_b1-signd_b1:0] bb1 [nb_in_reg:0];
  reg [width_c1-signd_c1:0] cc1 [nb_in_reg:0];
  reg [width_d1-signd_d1:0] dd1 [nb_in_reg:0];
  reg [sop_len-1:0] sop [nb_sop_reg:0];

  reg [width_e-signd_e:0] ee [n_inreg:0];
  reg                     accum [n_inreg:0];
  reg                     vl [n_inreg:0];

  genvar i;

  // make all inputs signed
  always @(*) aa0[nb_in_reg] = signd_a0 ? a0 : {1'b0, a0};
  always @(*) bb0[nb_in_reg] = signd_b0 ? b0 : {1'b0, b0};
  always @(*) cc0[nb_in_reg] = signd_c0 ? c0 : {1'b0, c0};
  generate if (width_d1>0 && width_d0>0) begin
    always @(*) dd0[nb_in_reg] = signd_d0 ? d0 : {1'b0, d0};
  end endgenerate
  always @(*) aa1[nb_in_reg] = signd_a1 ? a1 : {1'b0, a1};
  always @(*) bb1[nb_in_reg] = signd_b1 ? b1 : {1'b0, b1};
  always @(*) cc1[nb_in_reg] = signd_c1 ? c1 : {1'b0, c1};
  generate if (width_d1>0 && width_d0>0) begin
    always @(*) dd1[nb_in_reg] = signd_d1 ? d1 : {1'b0, d1};
  end endgenerate
  always @(*) ee[nb_in_reg] = signd_e ? e : {1'b0, e};
  always @(*) accum[n_inreg] = !load;
  always @(*) vl[n_inreg] = datavalid;

  // input registers
  generate if (n_inreg>0) begin
  for(i = n_inreg-1; i >= 0; i=i-1) begin:in_pipe_prod
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) aa0[i] <= aa0[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) aa1[i] <= aa1[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) bb0[i] <= bb0[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) bb1[i] <= bb1[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) cc0[i] <= cc0[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) cc1[i] <= cc1[i+1];//spyglass disable FlopEConst
      if (width_d0>0 && width_d1>0) begin
        always @(posedge(clk)) if (en == enable_active) dd0[i] <= dd0[i+1];//spyglass disable FlopEConst
        always @(posedge(clk)) if (en == enable_active) dd1[i] <= dd1[i+1];//spyglass disable FlopEConst
      end
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) aa0[i] <= aa0[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) aa1[i] <= aa1[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) bb0[i] <= bb0[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) bb1[i] <= bb1[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) cc0[i] <= cc0[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) cc1[i] <= cc1[i+1];//spyglass disable FlopEConst
      if (width_d0>0 && width_d1>0) begin
        always @(negedge(clk)) if (en == enable_active) dd0[i] <= dd0[i+1];//spyglass disable FlopEConst
        always @(negedge(clk)) if (en == enable_active) dd1[i] <= dd1[i+1];//spyglass disable FlopEConst
      end
    end
  end end endgenerate

  generate if (n_inreg>0) begin
  for(i = n_inreg-1; i >= 0; i=i-1) begin:in_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) accum[i] <= accum[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) vl[i] <= vl[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) accum[i] <= accum[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) vl[i] <= vl[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // perform products
  reg  [width_a0-signd_a0+1+width_a1-signd_a1+1-1:0] xa[nb_prod_reg:0];
  reg  [width_b0-signd_b0+1+width_b1-signd_b1+1-1:0] xb[nb_prod_reg:0];
  reg  [width_c0-signd_c0+1+width_c1-signd_c1+1-1:0] xc[nb_prod_reg:0];
  reg  [width_d0-signd_d0+1+width_d1-signd_d1+1-1:0] xd[nb_prod_reg:0];
  always @(*) xa[nb_prod_reg] = $signed(aa0[0]) * $signed(aa1[0]);
  always @(*) xb[nb_prod_reg] = $signed(bb0[0]) * $signed(bb1[0]);
  always @(*) xc[nb_prod_reg] = $signed(cc0[0]) * $signed(cc1[0]);
  generate if (nb_prod_reg>0) begin
  for(i = nb_prod_reg-1; i >= 0; i=i-1) begin:prod_pipe1
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) xa[i] <= xa[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) xb[i] <= xb[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) xc[i] <= xc[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) xa[i] <= xa[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) xb[i] <= xb[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) xc[i] <= xc[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  generate if (width_d0>0 && width_d1>0) begin:prod_pipe2
    always @(*) xd[nb_prod_reg] = $signed(dd0[0]) * $signed(dd1[0]);
    if (nb_prod_reg>0) begin
    for(i = nb_prod_reg-1; i >= 0; i=i-1) begin:prod_pipe3
      if (clock_edge == 1'b1) begin:pos
        always @(posedge(clk)) if (en == enable_active) xd[i] <= xd[i+1];//spyglass disable FlopEConst
      end else begin:neg
        always @(negedge(clk)) if (en == enable_active) xd[i] <= xd[i+1];//spyglass disable FlopEConst
      end
    end end
  end endgenerate


  generate
    if ( width_d0>0 && width_d1>0)       always @(*) sop[nb_sop_reg] = proda_pol*$signed(xa[0]) + prodb_pol*$signed(xb[0]) + prodc_pol*$signed(xc[0]) + prodd_pol*$signed(xd[0]);
    if ( width_d0==0 && width_d1==0) begin
      // Not supported by Vivado2020.2 : always @(*) sop[sumofprod_stages] = proda_pol*$signed(xa[0]) + prodb_pol*$signed(xb[0]) + prodc_pol*$signed(c1xc2[0]);
      if ( add_a==1 && add_b==1 && add_c==1) always @(*) sop[nb_sop_reg] = $signed(xa[0]) + $signed(xb[0]) + $signed(xc[0]);
      if ( add_a==1 && add_b==1 && add_c==0) always @(*) sop[nb_sop_reg] = $signed(xa[0]) + $signed(xb[0]) - $signed(xc[0]);
      if ( add_a==1 && add_b==0 && add_c==1) always @(*) sop[nb_sop_reg] = $signed(xa[0]) - $signed(xb[0]) + $signed(xc[0]);
      if ( add_a==1 && add_b==0 && add_c==0) always @(*) sop[nb_sop_reg] = $signed(xa[0]) - $signed(xb[0]) - $signed(xc[0]);
      if ( add_a==0 && add_b==1 && add_c==1) always @(*) sop[nb_sop_reg] = -$signed(xa[0]) + $signed(xb[0]) + $signed(xc[0]);
      if ( add_a==0 && add_b==1 && add_c==0) always @(*) sop[nb_sop_reg] = -$signed(xa[0]) + $signed(xb[0]) - $signed(xc[0]);
      if ( add_a==0 && add_b==0 && add_c==1) always @(*) sop[nb_sop_reg] = -$signed(xa[0]) - $signed(xb[0]) + $signed(xc[0]);
      if ( add_a==0 && add_b==0 && add_c==0) always @(*) sop[nb_sop_reg] = -$signed(xa[0]) - $signed(xb[0]) - $signed(xc[0]);
    end
  endgenerate
  generate if (nb_sop_reg>0) begin
  for(i = nb_sop_reg-1; i >= 0; i=i-1) begin:sop_pipe1
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) sop[i] <= sop[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) sop[i] <= sop[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg  [zz_len-1:0]  zz[out_stages-1:0];
  wire [zz_len-1:0]  z_or_e;
  assign z_or_e = accum[0] ? $signed(zz[out_stages-2]) : $signed(ee[0]);
  always @(*) zz[out_stages-1] = $signed(z_or_e) + $signed(sop[0]);

  // Output registers:
  generate if (out_stages>1) begin
  for(i = out_stages-2; i >= 0; i=i-1) begin:out_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active && (vl[0] || i != out_stages-2)) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active && (vl[0] || i != out_stages-2)) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // adjust output
  assign z = zz[0];

endmodule // mgc_mul4acc_pipe

//------> /cad/mentor/2024.2_1/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)
// suppress_sim_read_addr_range_errs:  0 - report errors  1 - suppress errors

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 ,
  parameter suppress_sim_read_addr_range_errs = 1 
  
)( clk,clken,d,q,radr,re,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input  re;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" , syn_ramstyle = "block" *)
  reg [data_width-1:0] mem [depth-1:0];
  integer j;
  initial for (j = 0; j < depth; j = j + 1) mem[j] = 0;
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr READ_ENABLE re
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg re_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
          re_reg <= re;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./PECore.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   code@iron-06
//  Generated date: Thu Jan 15 14:43:00 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_139_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_139_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_PECoreRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_PECoreRun_fsm (
  clk, rst, PECoreRun_wen, fsm_output
);
  input clk;
  input rst;
  input PECoreRun_wen;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for PECore_PECore_PECoreRun_PECoreRun_fsm_1
  parameter
    PECoreRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : PECore_PECore_PECoreRun_PECoreRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // PECoreRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= PECoreRun_rlp_C_0;
    end
    else if ( PECoreRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_staller
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_staller (
  clk, rst, PECoreRun_wen, PECoreRun_wten, act_port_Push_mioi_wen_comp, rva_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PECoreRun_wen;
  output PECoreRun_wten;
  input act_port_Push_mioi_wen_comp;
  input rva_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg PECoreRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign PECoreRun_wen = act_port_Push_mioi_wen_comp & rva_out_Push_mioi_wen_comp;
  assign PECoreRun_wten = PECoreRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECoreRun_wten_reg <= 1'b0;
    end
    else begin
      PECoreRun_wten_reg <= ~ PECoreRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_wait_dp (
  weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      ProductSum_for_acc_20_cmp_en, ProductSum_for_acc_19_cmp_en, PECoreRun_wen,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg,
      PECore_RunScale_if_for_4_mul_1_cmp_cgo, PECore_RunScale_if_for_4_mul_1_cmp_cgo_ir_unreg,
      PECore_RunScale_if_for_4_mul_1_cmp_en, ProductSum_for_acc_20_cmp_cgo, ProductSum_for_acc_20_cmp_cgo_ir_unreg,
      ProductSum_for_acc_19_cmp_cgo, ProductSum_for_acc_19_cmp_cgo_ir_unreg
);
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output ProductSum_for_acc_20_cmp_en;
  output ProductSum_for_acc_19_cmp_en;
  input PECoreRun_wen;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg;
  input PECore_RunScale_if_for_4_mul_1_cmp_cgo;
  input PECore_RunScale_if_for_4_mul_1_cmp_cgo_ir_unreg;
  output PECore_RunScale_if_for_4_mul_1_cmp_en;
  input ProductSum_for_acc_20_cmp_cgo;
  input ProductSum_for_acc_20_cmp_cgo_ir_unreg;
  input ProductSum_for_acc_19_cmp_cgo;
  input ProductSum_for_acc_19_cmp_cgo_ir_unreg;



  // Interconnect Declarations for Component Instantiations 
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg);
  assign PECore_RunScale_if_for_4_mul_1_cmp_en = PECoreRun_wen & (PECore_RunScale_if_for_4_mul_1_cmp_cgo
      | PECore_RunScale_if_for_4_mul_1_cmp_cgo_ir_unreg);
  assign ProductSum_for_acc_20_cmp_en = ~(PECoreRun_wen & (ProductSum_for_acc_20_cmp_cgo
      | ProductSum_for_acc_20_cmp_cgo_ir_unreg));
  assign ProductSum_for_acc_19_cmp_en = ~(PECoreRun_wen & (ProductSum_for_acc_19_cmp_cgo
      | ProductSum_for_acc_19_cmp_cgo_ir_unreg));
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  PECoreRun_wen, rva_out_Push_mioi_oswt, rva_out_Push_mioi_biwt, rva_out_Push_mioi_bdwt,
      rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & PECoreRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt)
      & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & rva_out_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt,
      start_PopNB_mioi_biwt_pff, start_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_biwt_pff;
  input start_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & PECoreRun_wen;
  assign start_PopNB_mioi_biwt = (~ PECoreRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_biwt_pff = PECoreRun_wen & start_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp (
  clk, rst, act_port_Push_mioi_oswt, act_port_Push_mioi_wen_comp, act_port_Push_mioi_biwt,
      act_port_Push_mioi_bdwt, act_port_Push_mioi_bcwt
);
  input clk;
  input rst;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input act_port_Push_mioi_biwt;
  input act_port_Push_mioi_bdwt;
  output act_port_Push_mioi_bcwt;
  reg act_port_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_wen_comp = (~ act_port_Push_mioi_oswt) | act_port_Push_mioi_biwt
      | act_port_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_Push_mioi_bcwt <= ~((~(act_port_Push_mioi_bcwt | act_port_Push_mioi_biwt))
          | act_port_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl (
  PECoreRun_wen, act_port_Push_mioi_oswt, act_port_Push_mioi_biwt, act_port_Push_mioi_bdwt,
      act_port_Push_mioi_bcwt, act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      act_port_Push_mioi_ccs_ccore_done_sync_vld, act_port_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_biwt;
  output act_port_Push_mioi_bdwt;
  input act_port_Push_mioi_bcwt;
  output act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input act_port_Push_mioi_ccs_ccore_done_sync_vld;
  input act_port_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_bdwt = act_port_Push_mioi_oswt & PECoreRun_wen;
  assign act_port_Push_mioi_biwt = act_port_Push_mioi_oswt & (~ act_port_Push_mioi_bcwt)
      & act_port_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & act_port_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
    (
  clk, rst, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt,
      input_port_PopNB_mioi_return_rsc_z_mxwt, input_port_PopNB_mioi_biwt, input_port_PopNB_mioi_bdwt,
      input_port_PopNB_mioi_data_data_data_rsc_z, input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_biwt;
  input input_port_PopNB_mioi_bdwt;
  input [127:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  input [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  input input_port_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg input_port_PopNB_mioi_bcwt;
  reg [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_bfwt;
  reg [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt;
  reg input_port_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_data_data_data_rsc_z_mxwt = MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z,
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt = MUX_v_8_2_2(input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z,
      input_port_PopNB_mioi_return_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      input_port_PopNB_mioi_bcwt <= ~((~(input_port_PopNB_mioi_bcwt | input_port_PopNB_mioi_biwt))
          | input_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= 8'b00000000;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( input_port_PopNB_mioi_biwt ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= input_port_PopNB_mioi_data_data_data_rsc_z;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= input_port_PopNB_mioi_data_logical_addr_rsc_z;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= input_port_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
    (
  PECoreRun_wen, PECoreRun_wten, input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_biwt,
      input_port_PopNB_mioi_bdwt, input_port_PopNB_mioi_biwt_pff, input_port_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output input_port_PopNB_mioi_biwt;
  output input_port_PopNB_mioi_bdwt;
  output input_port_PopNB_mioi_biwt_pff;
  input input_port_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_bdwt = input_port_PopNB_mioi_oswt & PECoreRun_wen;
  assign input_port_PopNB_mioi_biwt = (~ PECoreRun_wten) & input_port_PopNB_mioi_oswt;
  assign input_port_PopNB_mioi_biwt_pff = PECoreRun_wen & input_port_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [127:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  reg [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_128_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_20_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4, rva_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= 20'b00000000000000000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & PECoreRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ PECoreRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = PECoreRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, PECoreRun_wen, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_PECoreRun, rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [127:0] rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_oswt_pff(rva_out_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi (
  clk, rst, start_vld, start_rdy, start_dat, PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_vld(start_vld),
      .this_rdy(start_rdy),
      .this_dat(start_dat),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_biwt_pff(start_PopNB_mioi_biwt_iff),
      .start_PopNB_mioi_oswt_pff(start_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi (
  clk, rst, act_port_vld, act_port_rdy, act_port_dat, PECoreRun_wen, act_port_Push_mioi_oswt,
      act_port_Push_mioi_wen_comp, act_port_Push_mioi_m_data_rsc_dat_PECoreRun, act_port_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input [255:0] act_port_Push_mioi_m_data_rsc_dat_PECoreRun;
  input act_port_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_port_Push_mioi_biwt;
  wire act_port_Push_mioi_bdwt;
  wire act_port_Push_mioi_bcwt;
  wire act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire act_port_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push  act_port_Push_mioi
      (
      .this_vld(act_port_vld),
      .this_rdy(act_port_rdy),
      .this_dat(act_port_dat),
      .m_data_rsc_dat(act_port_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt),
      .act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .act_port_Push_mioi_ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .act_port_Push_mioi_oswt_pff(act_port_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi (
  clk, rst, input_port_vld, input_port_rdy, input_port_dat, PECoreRun_wen, PECoreRun_wten,
      input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt, input_port_PopNB_mioi_return_rsc_z_mxwt,
      input_port_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input input_port_vld;
  output input_port_rdy;
  input [137:0] input_port_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_port_PopNB_mioi_biwt;
  wire input_port_PopNB_mioi_bdwt;
  wire [127:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  wire input_port_PopNB_mioi_return_rsc_z;
  wire input_port_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB  input_port_PopNB_mioi
      (
      .this_vld(input_port_vld),
      .this_rdy(input_port_rdy),
      .this_dat(input_port_dat),
      .data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .return_rsc_z(input_port_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(input_port_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(input_port_PopNB_mioi_oswt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_biwt_pff(input_port_PopNB_mioi_biwt_iff),
      .input_port_PopNB_mioi_oswt_pff(input_port_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .input_port_PopNB_mioi_return_rsc_z(input_port_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt,
      rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG, weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d, ProductSum_for_acc_20_cmp_a,
      ProductSum_for_acc_20_cmp_load, ProductSum_for_acc_20_cmp_en, ProductSum_for_acc_20_cmp_z,
      ProductSum_for_acc_19_cmp_a0, ProductSum_for_acc_19_cmp_b0, ProductSum_for_acc_19_cmp_c0,
      ProductSum_for_acc_19_cmp_en, ProductSum_for_acc_19_cmp_z, ProductSum_for_acc_18_cmp_a0,
      ProductSum_for_acc_18_cmp_b0, ProductSum_for_acc_18_cmp_c0, ProductSum_for_acc_18_cmp_z,
      ProductSum_for_acc_17_cmp_a0, ProductSum_for_acc_17_cmp_b0, ProductSum_for_acc_17_cmp_c0,
      ProductSum_for_acc_17_cmp_z, ProductSum_for_acc_16_cmp_a0, ProductSum_for_acc_16_cmp_b0,
      ProductSum_for_acc_16_cmp_c0, ProductSum_for_acc_16_cmp_z, ProductSum_for_acc_15_cmp_a0,
      ProductSum_for_acc_15_cmp_b0, ProductSum_for_acc_15_cmp_c0, ProductSum_for_acc_15_cmp_z,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_a, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_load,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_z, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_a0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_b0, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_c0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_z, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_b0, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_c0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_b0, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_c0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_a,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_load, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_z,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_a0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_b0,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_c0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_b0,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_c0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_b0,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_c0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_a, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_z,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_a0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_b0,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_c0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_b0,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_c0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_b0,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_c0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_a, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_load,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_z, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_a0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_b0, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_c0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_z, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_b0, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_c0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_b0, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_c0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_a,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_z, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_a0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_b0, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_c0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_z, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_b0, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_c0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b0, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_c0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_a,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_load, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_z,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_a0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_b0,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_c0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_b0,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_c0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_b0,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_c0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_a, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_load,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_z, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_a0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_b0, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_c0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_z, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_b0, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_c0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_b0, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_c0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z, ProductSum_for_acc_20_cmp_b_pff,
      ProductSum_for_acc_20_cmp_datavalid_pff, ProductSum_for_acc_19_cmp_a1_pff,
      ProductSum_for_acc_19_cmp_b1_pff, ProductSum_for_acc_19_cmp_c1_pff, ProductSum_for_acc_19_cmp_load_pff,
      ProductSum_for_acc_19_cmp_datavalid_pff, ProductSum_for_acc_18_cmp_a1_pff,
      ProductSum_for_acc_18_cmp_b1_pff, ProductSum_for_acc_18_cmp_c1_pff, ProductSum_for_acc_17_cmp_a1_pff,
      ProductSum_for_acc_17_cmp_b1_pff, ProductSum_for_acc_17_cmp_c1_pff, ProductSum_for_acc_16_cmp_a1_pff,
      ProductSum_for_acc_16_cmp_b1_pff, ProductSum_for_acc_16_cmp_c1_pff, ProductSum_for_acc_15_cmp_a1_pff,
      ProductSum_for_acc_15_cmp_b1_pff, ProductSum_for_acc_15_cmp_c1_pff, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_pff,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_pff, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_b_pff,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_pff, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_pff,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_pff, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_pff,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff, weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [137:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  output [7:0] ProductSum_for_acc_20_cmp_a;
  output ProductSum_for_acc_20_cmp_load;
  output ProductSum_for_acc_20_cmp_en;
  input [30:0] ProductSum_for_acc_20_cmp_z;
  output [7:0] ProductSum_for_acc_19_cmp_a0;
  output [7:0] ProductSum_for_acc_19_cmp_b0;
  output [7:0] ProductSum_for_acc_19_cmp_c0;
  output ProductSum_for_acc_19_cmp_en;
  input [30:0] ProductSum_for_acc_19_cmp_z;
  output [7:0] ProductSum_for_acc_18_cmp_a0;
  output [7:0] ProductSum_for_acc_18_cmp_b0;
  output [7:0] ProductSum_for_acc_18_cmp_c0;
  input [30:0] ProductSum_for_acc_18_cmp_z;
  output [7:0] ProductSum_for_acc_17_cmp_a0;
  output [7:0] ProductSum_for_acc_17_cmp_b0;
  output [7:0] ProductSum_for_acc_17_cmp_c0;
  input [30:0] ProductSum_for_acc_17_cmp_z;
  output [7:0] ProductSum_for_acc_16_cmp_a0;
  output [7:0] ProductSum_for_acc_16_cmp_b0;
  output [7:0] ProductSum_for_acc_16_cmp_c0;
  input [30:0] ProductSum_for_acc_16_cmp_z;
  output [7:0] ProductSum_for_acc_15_cmp_a0;
  output [7:0] ProductSum_for_acc_15_cmp_b0;
  output [7:0] ProductSum_for_acc_15_cmp_c0;
  input [30:0] ProductSum_for_acc_15_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_a;
  output PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_load;
  input [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_a;
  output PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_load;
  input [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_a;
  input [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_a;
  output PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_load;
  input [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_a;
  input [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_a;
  output PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_load;
  input [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_a;
  output PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_load;
  input [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] ProductSum_for_acc_20_cmp_b_pff;
  output ProductSum_for_acc_20_cmp_datavalid_pff;
  output [7:0] ProductSum_for_acc_19_cmp_a1_pff;
  output [7:0] ProductSum_for_acc_19_cmp_b1_pff;
  output [7:0] ProductSum_for_acc_19_cmp_c1_pff;
  output ProductSum_for_acc_19_cmp_load_pff;
  output ProductSum_for_acc_19_cmp_datavalid_pff;
  output [7:0] ProductSum_for_acc_18_cmp_a1_pff;
  output [7:0] ProductSum_for_acc_18_cmp_b1_pff;
  output [7:0] ProductSum_for_acc_18_cmp_c1_pff;
  output [7:0] ProductSum_for_acc_17_cmp_a1_pff;
  output [7:0] ProductSum_for_acc_17_cmp_b1_pff;
  output [7:0] ProductSum_for_acc_17_cmp_c1_pff;
  output [7:0] ProductSum_for_acc_16_cmp_a1_pff;
  output [7:0] ProductSum_for_acc_16_cmp_b1_pff;
  output [7:0] ProductSum_for_acc_16_cmp_c1_pff;
  output [7:0] ProductSum_for_acc_15_cmp_a1_pff;
  output [7:0] ProductSum_for_acc_15_cmp_b1_pff;
  output [7:0] ProductSum_for_acc_15_cmp_c1_pff;
  output PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_pff;
  output PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_pff;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_b_pff;
  output PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_pff;
  output PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_pff;
  output PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_pff;
  output PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_pff;
  output PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff;


  // Interconnect Declarations
  wire PECoreRun_wen;
  wire PECoreRun_wten;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  wire input_port_PopNB_mioi_return_rsc_z_mxwt;
  wire act_port_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire PECore_RunScale_if_for_4_mul_1_cmp_en;
  wire [38:0] PECore_RunScale_if_for_4_mul_1_cmp_z;
  wire [38:0] PECore_RunScale_if_for_4_mul_1_cmp_1_z;
  wire [38:0] PECore_RunScale_if_for_4_mul_1_cmp_2_z;
  wire [38:0] PECore_RunScale_if_for_4_mul_1_cmp_3_z;
  wire [38:0] PECore_RunScale_if_for_4_mul_1_cmp_4_z;
  wire [38:0] PECore_RunScale_if_for_4_mul_1_cmp_5_z;
  wire [38:0] PECore_RunScale_if_for_4_mul_1_cmp_6_z;
  wire [38:0] PECore_RunScale_if_for_4_mul_1_cmp_7_z;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
  wire fsm_output;
  wire pe_config_UpdateManagerCounter_if_if_unequal_tmp;
  wire [7:0] weight_mem_write_arbxbar_xbar_for_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp;
  wire while_mux_1443_tmp;
  wire while_mux_1442_tmp;
  wire while_mux_1441_tmp;
  wire while_mux_1440_tmp;
  wire while_mux_1439_tmp;
  wire while_mux_1438_tmp;
  wire while_mux_1437_tmp;
  wire while_mux_1436_tmp;
  wire while_mux_1435_tmp;
  wire while_mux_1434_tmp;
  wire while_mux_1433_tmp;
  wire while_mux_1432_tmp;
  wire while_mux_1431_tmp;
  wire while_mux_1430_tmp;
  wire while_mux_1427_tmp;
  wire while_mux_1426_tmp;
  wire while_mux_1425_tmp;
  wire while_mux_1424_tmp;
  wire while_mux_1422_tmp;
  wire while_mux_1421_tmp;
  wire while_mux_1420_tmp;
  wire while_mux_1408_tmp;
  wire while_mux_1407_tmp;
  wire while_mux_1406_tmp;
  wire while_mux_1405_tmp;
  wire while_mux_1403_tmp;
  wire while_mux_1401_tmp;
  wire while_mux_1400_tmp;
  wire while_mux_1399_tmp;
  wire while_mux_1398_tmp;
  wire while_mux_1396_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_123_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_111_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_99_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_91_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_75_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_60_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_56_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_34_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp;
  wire while_and_40_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  wire and_dcpl_6;
  wire and_dcpl_7;
  wire and_dcpl_8;
  wire and_dcpl_24;
  wire and_dcpl_29;
  wire or_tmp_8;
  wire and_dcpl_33;
  wire and_dcpl_35;
  wire or_tmp_14;
  wire or_tmp_15;
  wire and_dcpl_40;
  wire not_tmp_33;
  wire nor_tmp_2;
  wire and_dcpl_47;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire or_tmp_23;
  wire and_tmp_1;
  wire or_tmp_24;
  wire or_dcpl_12;
  wire and_dcpl_76;
  wire and_dcpl_82;
  wire and_dcpl_84;
  wire and_dcpl_86;
  wire and_dcpl_88;
  wire or_dcpl_41;
  wire and_dcpl_90;
  wire or_dcpl_48;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_96;
  wire and_dcpl_98;
  wire and_dcpl_155;
  wire and_dcpl_162;
  wire and_dcpl_171;
  wire and_dcpl_174;
  wire and_dcpl_175;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_181;
  wire and_dcpl_182;
  wire and_dcpl_185;
  wire and_dcpl_187;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_194;
  wire and_dcpl_196;
  wire and_dcpl_198;
  wire and_dcpl_200;
  wire and_dcpl_202;
  wire and_dcpl_205;
  wire and_dcpl_206;
  wire and_dcpl_209;
  wire and_dcpl_212;
  wire and_dcpl_213;
  wire or_dcpl_146;
  wire and_dcpl_214;
  wire and_dcpl_218;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire and_dcpl_222;
  wire and_dcpl_224;
  wire or_tmp_36;
  wire or_tmp_37;
  wire and_dcpl_248;
  wire mux_tmp_42;
  wire mux_tmp_43;
  wire mux_tmp_47;
  wire mux_tmp_49;
  wire and_dcpl_262;
  wire and_dcpl_263;
  wire and_dcpl_277;
  wire and_dcpl_284;
  wire and_dcpl_290;
  wire and_dcpl_314;
  wire and_dcpl_323;
  wire and_dcpl_352;
  wire and_dcpl_353;
  wire and_dcpl_356;
  wire and_dcpl_382;
  wire or_tmp_85;
  wire or_dcpl_216;
  wire and_dcpl_415;
  wire and_dcpl_419;
  wire and_dcpl_421;
  wire or_tmp_108;
  wire and_dcpl_434;
  wire and_dcpl_445;
  wire or_tmp_112;
  wire not_tmp_248;
  wire and_dcpl_464;
  wire mux_tmp_95;
  wire and_dcpl_477;
  wire and_dcpl_497;
  wire and_dcpl_507;
  wire and_dcpl_514;
  wire and_tmp_4;
  wire and_dcpl_516;
  wire and_tmp_5;
  wire and_tmp_6;
  wire and_tmp_7;
  wire mux_tmp_108;
  wire and_tmp_8;
  wire and_tmp_9;
  wire and_tmp_10;
  wire mux_tmp_118;
  wire and_tmp_11;
  wire and_dcpl_539;
  wire and_dcpl_541;
  wire and_dcpl_552;
  wire and_dcpl_553;
  wire or_dcpl_243;
  wire or_dcpl_249;
  wire or_dcpl_251;
  wire or_dcpl_252;
  wire or_dcpl_253;
  wire or_dcpl_255;
  wire and_dcpl_576;
  wire or_dcpl_258;
  wire and_dcpl_593;
  wire and_dcpl_598;
  wire and_dcpl_615;
  wire and_dcpl_619;
  wire or_dcpl_259;
  wire or_dcpl_270;
  wire or_dcpl_271;
  wire and_dcpl_631;
  wire and_dcpl_632;
  wire and_dcpl_633;
  wire and_dcpl_634;
  wire or_dcpl_305;
  wire and_dcpl_637;
  wire and_dcpl_638;
  wire or_dcpl_309;
  wire and_dcpl_658;
  wire and_dcpl_659;
  wire and_dcpl_663;
  wire or_tmp_187;
  wire mux_tmp_166;
  wire mux_tmp_167;
  wire mux_tmp_171;
  wire nand_tmp_8;
  wire mux_tmp_177;
  wire mux_tmp_178;
  wire mux_tmp_182;
  wire or_tmp_201;
  wire nor_tmp_65;
  wire mux_tmp_189;
  wire or_tmp_205;
  wire mux_tmp_190;
  wire nor_tmp_70;
  wire mux_tmp_192;
  wire mux_tmp_193;
  wire mux_tmp_194;
  wire mux_tmp_195;
  wire or_tmp_213;
  wire or_tmp_217;
  wire or_tmp_225;
  wire mux_tmp_209;
  wire or_tmp_232;
  wire and_dcpl_672;
  wire or_tmp_239;
  wire or_tmp_241;
  wire mux_tmp_220;
  wire mux_tmp_223;
  wire mux_tmp_226;
  wire or_tmp_246;
  wire or_tmp_251;
  wire or_tmp_254;
  wire mux_tmp_233;
  wire or_tmp_258;
  wire or_tmp_264;
  wire or_tmp_270;
  wire and_dcpl_675;
  wire or_tmp_279;
  wire or_tmp_284;
  wire nor_tmp_118;
  wire nor_tmp_121;
  wire mux_tmp_254;
  wire or_tmp_296;
  wire or_tmp_297;
  wire or_tmp_304;
  wire or_tmp_305;
  wire not_tmp_441;
  wire or_tmp_312;
  wire or_tmp_318;
  wire and_dcpl_678;
  wire nor_tmp_158;
  wire nor_tmp_159;
  wire or_dcpl_320;
  wire or_tmp_335;
  wire or_tmp_338;
  wire mux_tmp_290;
  wire or_tmp_341;
  wire or_tmp_345;
  wire or_tmp_346;
  wire and_dcpl_679;
  wire or_tmp_352;
  wire or_tmp_353;
  wire or_tmp_355;
  wire or_tmp_361;
  wire and_dcpl_680;
  wire or_tmp_369;
  wire mux_tmp_306;
  wire mux_tmp_307;
  wire mux_tmp_309;
  wire and_dcpl_684;
  wire or_tmp_377;
  wire or_tmp_379;
  wire and_dcpl_687;
  wire nor_tmp_195;
  wire or_tmp_381;
  wire or_tmp_382;
  wire nor_tmp_198;
  wire or_tmp_384;
  wire or_tmp_385;
  wire mux_tmp_321;
  wire mux_tmp_323;
  wire and_dcpl_688;
  wire and_dcpl_689;
  wire and_dcpl_695;
  wire nor_tmp_200;
  wire mux_tmp_330;
  wire or_tmp_397;
  wire mux_tmp_333;
  wire nor_tmp_209;
  wire or_tmp_399;
  wire or_tmp_400;
  wire or_tmp_401;
  wire mux_tmp_334;
  wire or_tmp_407;
  wire or_tmp_408;
  wire or_tmp_409;
  wire or_tmp_411;
  wire or_tmp_413;
  wire or_tmp_415;
  wire mux_tmp_338;
  wire or_tmp_418;
  wire or_tmp_419;
  wire mux_tmp_339;
  wire nand_tmp_17;
  wire and_dcpl_697;
  wire nor_tmp_224;
  wire or_tmp_436;
  wire mux_tmp_358;
  wire mux_tmp_359;
  wire mux_tmp_360;
  wire mux_tmp_363;
  wire nor_tmp_227;
  wire or_tmp_441;
  wire or_tmp_442;
  wire mux_tmp_364;
  wire mux_tmp_365;
  wire mux_tmp_366;
  wire or_tmp_447;
  wire or_tmp_450;
  wire mux_tmp_376;
  wire or_tmp_452;
  wire mux_tmp_377;
  wire or_tmp_460;
  wire not_tmp_470;
  wire or_tmp_467;
  wire or_tmp_473;
  wire and_dcpl_700;
  wire and_dcpl_704;
  wire and_dcpl_705;
  wire and_dcpl_708;
  wire or_dcpl_328;
  wire [3:0] pe_config_manager_counter_sva_mx1;
  wire [4:0] operator_4_false_acc_sdt_sva_1;
  wire [5:0] nl_operator_4_false_acc_sdt_sva_1;
  reg [3:0] pe_config_num_manager_sva;
  wire state_0_sva_mx1;
  wire while_if_and_tmp_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiWrite_switch_lp_nor_tmp_1;
  reg pe_config_is_valid_sva;
  reg pe_config_is_zero_first_sva;
  reg pe_manager_zero_active_sva;
  reg pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  reg pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  reg PECore_UpdateFSM_switch_lp_and_7_itm_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
  reg PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  reg [8:0] operator_8_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_8_false_acc_sdt_sva_1;
  wire PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  wire PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1;
  reg PECore_RunFSM_switch_lp_nor_tmp_1;
  reg [1:0] state_2_1_sva;
  reg state_0_sva;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  reg PECore_RunFSM_switch_lp_equal_tmp_1_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  reg weight_mem_run_3_for_land_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  reg input_read_req_valid_lpi_1_dfm_1_9;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
  reg rva_in_reg_rw_sva_9;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  wire PECore_UpdateFSM_switch_lp_equal_tmp_6;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  wire PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
  wire PECore_UpdateFSM_switch_lp_nor_tmp_1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
  wire [7:0] pe_config_input_counter_sva_mx1;
  wire [8:0] operator_16_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_16_false_acc_sdt_sva_1;
  reg [7:0] pe_manager_num_input_sva;
  reg [7:0] pe_config_num_output_sva;
  wire PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  wire PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0;
  reg PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
  wire weight_mem_run_3_for_land_lpi_1_dfm_1;
  wire weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  wire weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  wire weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_lpi_1_dfm_1_1;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_371_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1;
  wire weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1;
  reg rva_in_reg_rw_sva_5;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_127_sva_1;
  reg input_write_req_valid_lpi_1_dfm_1_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1;
  wire input_write_req_valid_lpi_1_dfm_5;
  wire input_mem_banks_write_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1;
  reg [14:0] pe_manager_base_input_sva;
  reg accum_vector_data_7_sva_1_load;
  reg accum_vector_data_6_sva_1_load;
  reg accum_vector_data_5_sva_1_load;
  reg accum_vector_data_4_sva_1_load;
  reg accum_vector_data_3_sva_1_load;
  reg accum_vector_data_2_sva_1_load;
  reg accum_vector_data_1_sva_1_load;
  reg accum_vector_data_0_sva_1_load;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_4;
  wire PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0;
  wire PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_mx0w0;
  reg rva_in_reg_rw_sva_st_1_9;
  reg while_stage_0_11;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
  reg input_read_req_valid_lpi_1_dfm_1_8;
  reg rva_in_reg_rw_sva_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  reg rva_in_reg_rw_sva_st_1_8;
  reg rva_in_reg_rw_sva_st_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  reg while_stage_0_10;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_8;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_1;
  reg while_stage_0_3;
  reg while_stage_0_4;
  reg while_stage_0_5;
  reg while_stage_0_6;
  reg while_stage_0_7;
  reg while_stage_0_8;
  reg while_stage_0_9;
  reg rva_in_reg_rw_sva_st_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  reg rva_in_reg_rw_sva_st_1_5;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
  reg ProductSum_for_asn_108_itm_3;
  reg ProductSum_for_asn_128_itm_3;
  reg ProductSum_for_asn_28_itm_3;
  reg ProductSum_for_asn_41_itm_3;
  reg ProductSum_for_asn_56_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
  reg ProductSum_for_asn_69_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3;
  reg PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  reg rva_in_reg_rw_sva_st_1_7;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_1;
  reg rva_in_reg_rw_sva_st_1_4;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_1_sva;
  reg rva_in_reg_rw_sva_st_7;
  reg input_read_req_valid_lpi_1_dfm_1_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
  reg rva_in_reg_rw_sva_7;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
  reg rva_in_reg_rw_sva_st_4;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
  reg rva_in_reg_rw_sva_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1;
  reg rva_in_reg_rw_sva_st_1_6;
  reg rva_in_reg_rw_sva_st_6;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
  reg input_read_req_valid_lpi_1_dfm_1_6;
  reg rva_in_reg_rw_sva_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5;
  reg rva_in_reg_rw_sva_3;
  reg accum_vector_operator_1_for_asn_73_itm_1;
  reg ProductSum_for_asn_56_itm_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
  reg [3:0] while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_9;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1;
  reg [1:0] state_2_1_sva_dfm_1;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_2;
  reg while_and_1263_itm_1;
  reg [7:0] weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_7_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_2_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_0_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_6_sva;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs;
  wire operator_7_false_1_operator_7_false_1_or_mdf_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_1_sva_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_3_2_0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_2_2_0;
  reg [14:0] weight_read_addrs_7_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_5_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_3_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_1_lpi_1_dfm_1;
  reg [14:0] pe_manager_base_weight_sva;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_2_2_0;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  wire [11:0] nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_2;
  wire [3:0] pe_manager_base_weight_sva_mx1_3_0;
  wire pe_manager_base_weight_sva_mx3_0;
  wire [14:0] pe_manager_base_weight_sva_mx2;
  reg [7:0] while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4;
  wire [7:0] input_write_addrs_lpi_1_dfm_2;
  wire PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
  wire Arbiter_8U_Roundrobin_pick_1_mux_133_mx1w1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_9_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_1_mux_63_mx1w1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_1_mux_62_mx1w1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1;
  wire while_and_221_rgt;
  wire while_and_225_rgt;
  wire while_and_229_rgt;
  wire while_and_233_rgt;
  wire while_and_237_rgt;
  wire while_and_241_rgt;
  wire while_and_245_rgt;
  wire while_and_249_rgt;
  wire while_and_253_rgt;
  wire while_and_257_rgt;
  wire while_and_261_rgt;
  wire while_and_265_rgt;
  wire while_and_269_rgt;
  wire while_and_273_rgt;
  wire while_and_277_rgt;
  wire while_and_281_rgt;
  wire while_and_285_rgt;
  wire while_and_289_rgt;
  wire while_and_293_rgt;
  wire while_and_297_rgt;
  wire while_and_301_rgt;
  wire while_and_305_rgt;
  wire while_and_309_rgt;
  wire while_and_313_rgt;
  wire while_and_317_rgt;
  wire while_and_321_rgt;
  wire while_and_325_rgt;
  wire while_and_329_rgt;
  wire while_and_333_rgt;
  wire while_and_337_rgt;
  wire while_and_341_rgt;
  wire while_and_345_rgt;
  wire while_and_349_rgt;
  wire while_and_353_rgt;
  wire while_and_357_rgt;
  wire while_and_361_rgt;
  wire while_and_365_rgt;
  wire while_and_369_rgt;
  wire while_and_373_rgt;
  wire while_and_377_rgt;
  wire while_and_381_rgt;
  wire while_and_385_rgt;
  wire while_and_389_rgt;
  wire while_and_393_rgt;
  wire while_and_397_rgt;
  wire while_and_401_rgt;
  wire while_and_405_rgt;
  wire while_and_409_rgt;
  wire while_and_413_rgt;
  wire while_and_417_rgt;
  wire while_and_421_rgt;
  wire while_and_425_rgt;
  wire while_and_429_rgt;
  wire while_and_433_rgt;
  wire while_and_437_rgt;
  wire while_and_441_rgt;
  wire while_and_445_rgt;
  wire while_and_449_rgt;
  wire while_and_453_rgt;
  wire while_and_457_rgt;
  wire while_and_461_rgt;
  wire while_and_465_rgt;
  wire while_and_469_rgt;
  wire while_and_473_rgt;
  wire while_and_477_rgt;
  wire while_and_481_rgt;
  wire while_and_485_rgt;
  wire while_and_489_rgt;
  wire while_and_493_rgt;
  wire while_and_497_rgt;
  wire while_and_501_rgt;
  wire while_and_505_rgt;
  wire while_and_509_rgt;
  wire while_and_513_rgt;
  wire while_and_517_rgt;
  wire while_and_521_rgt;
  wire while_and_525_rgt;
  wire while_and_529_rgt;
  wire while_and_533_rgt;
  wire while_and_537_rgt;
  wire while_and_541_rgt;
  wire while_and_545_rgt;
  wire while_and_549_rgt;
  wire while_and_553_rgt;
  wire while_and_557_rgt;
  wire while_and_561_rgt;
  wire while_and_565_rgt;
  wire while_and_569_rgt;
  wire while_and_573_rgt;
  wire while_and_577_rgt;
  wire while_and_581_rgt;
  wire while_and_585_rgt;
  wire while_and_589_rgt;
  wire while_and_593_rgt;
  wire while_and_597_rgt;
  wire while_and_601_rgt;
  wire while_and_605_rgt;
  wire while_and_609_rgt;
  wire while_and_613_rgt;
  wire while_and_617_rgt;
  wire while_and_621_rgt;
  wire while_and_625_rgt;
  wire while_and_629_rgt;
  wire while_and_633_rgt;
  wire while_and_637_rgt;
  wire while_and_641_rgt;
  wire while_and_645_rgt;
  wire while_and_649_rgt;
  wire while_and_653_rgt;
  wire while_and_657_rgt;
  wire while_and_661_rgt;
  wire while_and_665_rgt;
  wire while_and_669_rgt;
  wire while_and_673_rgt;
  wire while_and_677_rgt;
  wire while_and_681_rgt;
  wire while_and_685_rgt;
  wire while_and_689_rgt;
  wire while_and_693_rgt;
  wire while_and_697_rgt;
  wire while_and_701_rgt;
  wire while_and_705_rgt;
  wire while_and_709_rgt;
  wire while_and_713_rgt;
  wire while_and_717_rgt;
  wire while_and_721_rgt;
  wire while_and_725_rgt;
  wire while_and_729_rgt;
  wire while_and_733_rgt;
  wire while_and_737_rgt;
  wire while_and_741_rgt;
  wire while_and_745_rgt;
  wire while_and_749_rgt;
  wire while_and_753_rgt;
  wire while_and_757_rgt;
  wire while_and_761_rgt;
  wire while_and_765_rgt;
  wire while_and_769_rgt;
  wire while_and_773_rgt;
  wire while_and_777_rgt;
  wire while_and_781_rgt;
  wire while_and_785_rgt;
  wire while_and_789_rgt;
  wire while_and_793_rgt;
  wire while_and_797_rgt;
  wire while_and_801_rgt;
  wire while_and_805_rgt;
  wire while_and_809_rgt;
  wire while_and_813_rgt;
  wire while_and_817_rgt;
  wire while_and_821_rgt;
  wire while_and_825_rgt;
  wire while_and_829_rgt;
  wire while_and_833_rgt;
  wire while_and_837_rgt;
  wire while_and_841_rgt;
  wire while_and_845_rgt;
  wire while_and_849_rgt;
  wire while_and_853_rgt;
  wire while_and_857_rgt;
  wire while_and_861_rgt;
  wire while_and_865_rgt;
  wire while_and_869_rgt;
  wire while_and_873_rgt;
  wire while_and_877_rgt;
  wire while_and_881_rgt;
  wire while_and_885_rgt;
  wire while_and_889_rgt;
  wire while_and_893_rgt;
  wire while_and_897_rgt;
  wire while_and_901_rgt;
  wire while_and_905_rgt;
  wire while_and_909_rgt;
  wire while_and_913_rgt;
  wire while_and_917_rgt;
  wire while_and_921_rgt;
  wire while_and_925_rgt;
  wire while_and_929_rgt;
  wire while_and_933_rgt;
  wire while_and_937_rgt;
  wire while_and_941_rgt;
  wire while_and_945_rgt;
  wire while_and_949_rgt;
  wire while_and_953_rgt;
  wire while_and_957_rgt;
  wire while_and_961_rgt;
  wire while_and_965_rgt;
  wire while_and_969_rgt;
  wire while_and_973_rgt;
  wire while_and_977_rgt;
  wire while_and_981_rgt;
  wire while_and_985_rgt;
  wire while_and_989_rgt;
  wire while_and_993_rgt;
  wire while_and_997_rgt;
  wire while_and_1001_rgt;
  wire while_and_1005_rgt;
  wire while_and_1009_rgt;
  wire while_and_1013_rgt;
  wire while_and_1017_rgt;
  wire while_and_1021_rgt;
  wire while_and_1025_rgt;
  wire while_and_1029_rgt;
  wire while_and_1033_rgt;
  wire while_and_1037_rgt;
  wire while_and_1041_rgt;
  wire while_and_1045_rgt;
  wire while_and_1049_rgt;
  wire while_and_1053_rgt;
  wire while_and_1057_rgt;
  wire while_and_1061_rgt;
  wire while_and_1065_rgt;
  wire while_and_1069_rgt;
  wire while_and_1073_rgt;
  wire while_and_1077_rgt;
  wire while_and_1081_rgt;
  wire while_and_1085_rgt;
  wire while_and_1089_rgt;
  wire while_and_1093_rgt;
  wire while_and_1097_rgt;
  wire while_and_1101_rgt;
  wire while_and_1105_rgt;
  wire while_and_1109_rgt;
  wire while_and_1113_rgt;
  wire while_and_1117_rgt;
  wire while_and_1121_rgt;
  wire while_and_1125_rgt;
  wire while_and_1129_rgt;
  wire while_and_1133_rgt;
  wire while_and_1137_rgt;
  wire while_and_1141_rgt;
  wire while_and_1145_rgt;
  wire while_and_1149_rgt;
  wire while_and_1153_rgt;
  wire while_and_1157_rgt;
  wire while_and_1161_rgt;
  wire while_and_1165_rgt;
  wire while_and_1169_rgt;
  wire while_and_1173_rgt;
  wire while_and_1177_rgt;
  wire while_and_1181_rgt;
  wire while_and_1185_rgt;
  wire while_and_1189_rgt;
  wire while_and_1193_rgt;
  wire while_and_1197_rgt;
  wire while_and_1201_rgt;
  wire while_and_1205_rgt;
  wire while_and_1209_rgt;
  wire while_and_1213_rgt;
  wire while_and_1217_rgt;
  wire while_and_1221_rgt;
  wire while_and_1225_rgt;
  wire while_and_1229_rgt;
  wire while_and_1233_rgt;
  wire while_and_1237_rgt;
  wire while_and_1241_rgt;
  wire weight_mem_banks_read_1_for_mux_cse;
  wire weight_mem_banks_read_1_for_mux_1_cse;
  wire weight_mem_banks_read_1_for_mux_4_cse;
  wire weight_mem_banks_read_1_for_mux_5_cse;
  wire weight_mem_banks_read_1_for_mux_8_cse;
  wire weight_mem_banks_read_1_for_mux_9_cse;
  wire weight_mem_banks_read_1_for_mux_12_cse;
  wire weight_mem_banks_read_1_for_mux_13_cse;
  wire weight_mem_banks_read_1_for_mux_16_cse;
  wire weight_mem_banks_read_1_for_mux_17_cse;
  wire weight_mem_banks_read_1_for_mux_20_cse;
  wire weight_mem_banks_read_1_for_mux_21_cse;
  wire weight_mem_banks_read_1_for_mux_24_cse;
  wire weight_mem_banks_read_1_for_mux_25_cse;
  wire weight_mem_banks_read_1_for_mux_28_cse;
  wire weight_mem_banks_read_1_for_mux_29_cse;
  wire weight_mem_banks_write_if_for_if_mux_8_cse;
  wire weight_mem_banks_write_if_for_if_mux_9_cse;
  wire weight_mem_banks_read_for_mux_cse;
  wire weight_mem_banks_read_for_mux_1_cse;
  wire weight_mem_banks_write_if_for_if_mux_12_cse;
  wire weight_mem_banks_write_if_for_if_mux_13_cse;
  wire weight_mem_banks_read_for_mux_4_cse;
  wire weight_mem_banks_read_for_mux_5_cse;
  wire weight_mem_banks_write_if_for_if_mux_16_cse;
  wire weight_mem_banks_write_if_for_if_mux_17_cse;
  wire weight_mem_banks_read_for_mux_8_cse;
  wire weight_mem_banks_read_for_mux_9_cse;
  wire weight_mem_banks_write_if_for_if_mux_20_cse;
  wire weight_mem_banks_write_if_for_if_mux_21_cse;
  wire weight_mem_banks_read_for_mux_12_cse;
  wire weight_mem_banks_read_for_mux_13_cse;
  wire weight_mem_banks_write_if_for_if_mux_24_cse;
  wire weight_mem_banks_write_if_for_if_mux_25_cse;
  wire weight_mem_banks_read_for_mux_16_cse;
  wire weight_mem_banks_read_for_mux_17_cse;
  wire weight_mem_banks_write_if_for_if_mux_28_cse;
  wire weight_mem_banks_write_if_for_if_mux_29_cse;
  wire weight_mem_banks_read_for_mux_20_cse;
  wire weight_mem_banks_read_for_mux_21_cse;
  wire weight_mem_banks_write_if_for_if_mux_32_cse;
  wire weight_mem_banks_write_if_for_if_mux_33_cse;
  wire weight_mem_banks_read_for_mux_24_cse;
  wire weight_mem_banks_read_for_mux_25_cse;
  wire weight_mem_banks_write_if_for_if_mux_36_cse;
  wire weight_mem_banks_write_if_for_if_mux_37_cse;
  wire weight_mem_banks_read_for_mux_28_cse;
  wire weight_mem_banks_read_for_mux_29_cse;
  wire input_mem_banks_write_1_if_for_if_mux_cse;
  wire input_mem_banks_write_1_if_for_if_mux_1_cse;
  wire input_mem_banks_read_1_for_mux_cse;
  wire input_mem_banks_read_1_for_mux_1_cse;
  wire input_mem_banks_write_if_for_if_mux_cse;
  wire input_mem_banks_write_if_for_if_mux_1_cse;
  wire input_mem_banks_read_for_mux_cse;
  wire input_mem_banks_read_for_mux_1_cse;
  reg reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_cgo_ir_cse;
  reg reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_cgo_ir_cse;
  reg reg_PECore_RunScale_if_for_4_mul_1_cmp_cgo_ir_7_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_act_port_Push_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire rva_out_reg_data_and_cse;
  wire weight_port_read_out_data_and_cse;
  wire weight_port_read_out_data_and_16_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_cse;
  reg reg_rva_in_reg_rw_sva_st_1_1_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_or_2_cse;
  reg [2:0] reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse;
  reg reg_weight_mem_run_3_for_5_and_16_itm_1_cse;
  reg reg_weight_mem_run_3_for_5_and_14_itm_1_cse;
  wire operator_15_false_1_and_cse;
  wire pe_config_num_manager_and_cse;
  wire PECore_DecodeAxiWrite_switch_lp_and_cse;
  wire or_260_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2_cse;
  reg reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse;
  wire and_724_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
  wire pe_manager_num_input_and_cse;
  wire or_407_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_52_cse;
  wire Arbiter_8U_Roundrobin_pick_and_42_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_40_cse;
  wire Arbiter_8U_Roundrobin_pick_and_36_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_20_cse;
  wire Arbiter_8U_Roundrobin_pick_and_26_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_14_cse;
  wire Arbiter_8U_Roundrobin_pick_and_23_cse;
  wire Arbiter_8U_Roundrobin_pick_or_2_cse;
  wire Arbiter_8U_Roundrobin_pick_and_5_cse;
  wire [1:0] state_mux_1_cse;
  wire nor_384_cse;
  wire and_315_cse;
  wire nand_41_cse;
  wire nor_375_cse;
  wire and_747_cse;
  wire and_749_cse;
  wire or_222_cse;
  wire and_545_cse;
  wire and_549_cse;
  wire and_745_cse;
  wire or_237_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse;
  wire and_743_cse;
  wire and_742_cse;
  wire and_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_3_or_cse;
  wire nor_374_cse;
  wire or_113_cse;
  wire or_106_cse;
  wire or_92_cse;
  wire or_85_cse;
  wire and_754_cse;
  wire while_and_1243_cse;
  wire while_while_nor_259_cse;
  wire nor_310_cse;
  wire nor_285_cse;
  wire nor_286_cse;
  wire nor_290_cse;
  wire nor_294_cse;
  wire nor_297_cse;
  wire and_135_cse;
  wire nor_302_cse;
  wire nor_308_cse;
  wire nor_309_cse;
  wire nor_306_cse;
  wire nor_307_cse;
  wire nand_34_cse;
  wire nor_352_cse;
  wire while_and_39_cse;
  wire and_968_cse;
  wire or_516_cse;
  wire and_772_cse;
  wire and_771_cse;
  wire and_763_cse;
  wire and_778_cse;
  wire and_777_cse;
  wire and_776_cse;
  wire and_765_cse;
  wire and_781_cse;
  wire and_799_cse;
  wire and_805_cse;
  wire and_801_cse;
  wire and_809_cse;
  wire and_814_cse;
  wire and_804_cse;
  wire and_818_cse;
  wire and_808_cse;
  wire and_806_cse;
  wire and_810_cse;
  wire and_972_cse;
  wire and_976_cse;
  wire and_838_cse;
  wire and_975_cse;
  wire and_836_cse;
  wire and_971_cse;
  wire and_969_cse;
  wire and_970_cse;
  wire and_851_cse;
  wire and_973_cse;
  wire and_974_cse;
  wire and_849_cse;
  wire and_871_cse;
  wire and_872_cse;
  wire and_869_cse;
  wire and_870_cse;
  wire and_874_cse;
  wire and_878_cse;
  wire and_879_cse;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse;
  wire and_736_cse;
  wire and_907_cse;
  wire and_909_cse;
  wire and_738_cse;
  wire and_744_cse;
  wire nand_66_cse;
  wire and_908_cse;
  wire and_979_cse;
  wire and_936_cse;
  wire and_978_cse;
  wire and_977_cse;
  wire and_981_cse;
  wire and_980_cse;
  wire and_947_cse;
  wire and_941_cse;
  wire and_951_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1;
  reg accum_vector_operator_1_for_asn_73_itm_2;
  reg accum_vector_operator_1_for_asn_28_itm_2;
  reg accum_vector_operator_1_for_asn_43_itm_2;
  wire while_if_and_2_m1c;
  wire weight_mem_run_3_for_5_and_159_cse;
  wire weight_mem_run_3_for_5_and_161_cse;
  wire PECore_DecodeAxiRead_switch_lp_nor_2_cse;
  wire pe_config_is_valid_and_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_cse;
  wire Arbiter_8U_Roundrobin_pick_and_44_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_65_cse;
  wire Arbiter_8U_Roundrobin_pick_and_56_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_74_cse;
  wire Arbiter_8U_Roundrobin_pick_and_61_cse;
  wire pe_config_input_counter_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse;
  wire and_572_cse;
  wire while_and_4_cse;
  wire and_156_cse;
  wire and_107_cse;
  wire and_114_cse;
  wire and_121_cse;
  wire and_142_cse;
  wire or_614_cse;
  wire or_616_cse;
  wire or_659_cse;
  wire or_660_cse;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1;
  wire PECore_DecodeAxiWrite_switch_lp_or_5_cse_1;
  wire weight_mem_run_3_for_5_and_cse;
  wire weight_mem_run_3_for_5_and_173_cse;
  wire weight_mem_run_3_for_5_and_174_cse;
  wire weight_mem_run_3_for_5_and_176_cse;
  wire weight_mem_run_3_for_5_and_178_cse;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2_cse;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0;
  wire weight_mem_run_3_for_5_and_179_cse;
  wire and_543_rmff;
  wire and_540_rmff;
  wire and_537_rmff;
  wire and_534_rmff;
  wire and_531_rmff;
  wire and_527_rmff;
  wire and_523_rmff;
  wire and_520_rmff;
  wire and_516_rmff;
  wire and_514_rmff;
  wire and_511_rmff;
  wire and_547_rmff;
  reg [30:0] accum_vector_data_3_sva;
  reg [30:0] accum_vector_data_7_sva;
  reg [30:0] accum_vector_data_0_sva;
  reg [30:0] accum_vector_data_6_sva;
  reg [30:0] accum_vector_data_1_sva;
  reg [30:0] accum_vector_data_5_sva;
  reg [30:0] accum_vector_data_2_sva;
  reg [30:0] accum_vector_data_4_sva;
  reg [7:0] pe_config_output_counter_sva;
  reg [7:0] pe_config_input_counter_sva;
  reg [7:0] rva_out_reg_data_95_88_sva_dfm_4_4;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4_4;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4_4;
  reg rva_out_reg_data_63_sva_dfm_4_4;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_4;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4_4;
  reg rva_out_reg_data_47_sva_dfm_4_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_4;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_4;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1;
  reg [27:0] act_port_reg_data_251_224_sva;
  reg [27:0] act_port_reg_data_219_192_sva;
  reg [27:0] act_port_reg_data_187_160_sva;
  reg [27:0] act_port_reg_data_155_128_sva;
  reg [27:0] act_port_reg_data_123_96_sva;
  reg [27:0] act_port_reg_data_91_64_sva;
  reg [27:0] act_port_reg_data_59_32_sva;
  reg [27:0] act_port_reg_data_27_0_sva;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_4;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0;
  reg weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
  reg [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1;
  reg [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1;
  reg [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1;
  reg weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
  wire [7:0] weight_port_read_out_data_7_1_sva_dfm_2;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
  reg ProductSum_for_asn_28_itm_5;
  reg [7:0] weight_port_read_out_data_7_2_sva_dfm_1;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_5;
  reg [7:0] weight_port_read_out_data_7_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_0_sva_dfm_1;
  reg ProductSum_for_asn_26_itm_6;
  reg [7:0] weight_port_read_out_data_7_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_8_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_9_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_13_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_10_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_11_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_15_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_12_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg ProductSum_for_asn_41_itm_5;
  reg [7:0] weight_mem_run_3_for_5_mux_98_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_99_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_96_itm_1;
  reg ProductSum_for_asn_40_itm_6;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4_1;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4_1;
  reg [7:0] rva_out_reg_data_95_88_sva_dfm_4_1;
  reg [7:0] weight_port_read_out_data_5_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg ProductSum_for_asn_56_itm_5;
  reg [7:0] weight_mem_run_3_for_5_mux_82_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_83_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_80_itm_1;
  reg ProductSum_for_asn_55_itm_6;
  reg [7:0] weight_mem_run_3_for_5_mux_87_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_84_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_85_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_88_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_89_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_86_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_93_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_90_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_91_itm_1;
  reg [7:0] weight_port_read_out_data_5_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_15_sva_dfm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_92_itm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg [7:0] weight_port_read_out_data_4_1_sva_dfm_1;
  reg ProductSum_for_asn_69_itm_6;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  reg [7:0] weight_port_read_out_data_4_2_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  reg [7:0] weight_port_read_out_data_4_3_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  reg [7:0] weight_port_read_out_data_4_0_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  reg [7:0] weight_port_read_out_data_4_7_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  reg [7:0] weight_port_read_out_data_4_4_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  reg [7:0] weight_port_read_out_data_4_5_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  reg [7:0] weight_port_read_out_data_4_8_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  reg [7:0] weight_port_read_out_data_4_9_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  reg [7:0] weight_port_read_out_data_4_6_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  reg [7:0] weight_port_read_out_data_4_13_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  reg [7:0] weight_port_read_out_data_4_10_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  reg [7:0] weight_port_read_out_data_4_11_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  reg [7:0] weight_port_read_out_data_4_14_sva_dfm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_79_itm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
  reg [7:0] weight_port_read_out_data_4_12_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg ProductSum_for_asn_82_itm_5;
  reg [7:0] weight_mem_run_3_for_5_mux_50_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_51_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_48_itm_1;
  reg ProductSum_for_asn_81_itm_6;
  reg [7:0] weight_mem_run_3_for_5_mux_55_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_52_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_53_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_56_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_57_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_54_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_61_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_58_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_59_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_62_itm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
  reg [7:0] weight_port_read_out_data_3_15_sva_dfm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_60_itm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg [7:0] weight_port_read_out_data_2_1_sva_dfm_1;
  reg ProductSum_for_asn_95_itm_6;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  reg [7:0] weight_port_read_out_data_2_2_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  reg [7:0] weight_port_read_out_data_2_3_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  reg [7:0] weight_port_read_out_data_2_0_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  reg [7:0] weight_port_read_out_data_2_7_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  reg [7:0] weight_port_read_out_data_2_4_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  reg [7:0] weight_port_read_out_data_2_5_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  reg [7:0] weight_port_read_out_data_2_8_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  reg [7:0] weight_port_read_out_data_2_9_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  reg [7:0] weight_port_read_out_data_2_6_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  reg [7:0] weight_port_read_out_data_2_13_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  reg [7:0] weight_port_read_out_data_2_10_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  reg [7:0] weight_port_read_out_data_2_11_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  reg [7:0] weight_port_read_out_data_2_14_sva_dfm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_47_itm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
  reg [7:0] weight_port_read_out_data_2_12_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg ProductSum_for_asn_108_itm_5;
  reg [7:0] weight_mem_run_3_for_5_mux_18_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_19_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_16_itm_1;
  reg ProductSum_for_asn_107_itm_6;
  reg [7:0] weight_mem_run_3_for_5_mux_23_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_20_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_21_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_24_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_25_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_22_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_29_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_26_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_27_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_30_itm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
  reg [7:0] weight_port_read_out_data_1_15_sva_dfm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_28_itm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg ProductSum_for_asn_128_itm_5;
  reg ProductSum_for_asn_126_itm_6;
  reg [7:0] weight_port_read_out_data_0_7_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_0_5_sva_dfm_1_1;
  reg [7:0] weight_mem_run_3_for_5_mux_8_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_9_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_6_itm_1;
  reg [7:0] weight_write_data_data_0_15_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_14_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_13_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_12_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_11_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_10_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_9_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_8_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
  reg [14:0] weight_write_addrs_lpi_1_dfm_1_2;
  reg [7:0] weight_write_data_data_0_15_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_14_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_13_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_12_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_11_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_10_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_9_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_8_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_3_2;
  reg [11:0] weight_write_addrs_lpi_1_dfm_1_3_14_3;
  wire and_dcpl;
  wire and_dcpl_709;
  wire or_dcpl;
  wire or_dcpl_329;
  wire or_dcpl_331;
  wire or_dcpl_333;
  wire or_dcpl_334;
  wire and_dcpl_721;
  wire and_651_ssc;
  wire and_652_ssc;
  wire and_653_ssc;
  wire and_655_ssc;
  wire and_658_ssc;
  wire and_661_ssc;
  reg [127:0] input_mem_banks_read_read_data_lpi_1_dfm_1_4;
  reg [127:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1;
  wire [127:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0;
  wire [119:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_5;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1;
  wire or_847_tmp;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_4;
  wire and_1006_cse;
  wire and_1007_cse;
  wire and_1008_cse;
  wire and_1009_cse;
  wire and_1010_cse;
  wire and_1011_cse;
  wire nor_506_cse;
  wire and_1030_cse;
  wire and_1031_cse;
  wire and_1032_cse;
  wire and_1023_cse;
  wire and_1024_cse;
  wire and_1025_cse;
  wire and_1026_cse;
  wire and_1027_cse;
  wire nor_508_cse;
  wire [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm;
  wire [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm;
  wire [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm;
  wire mux_15_itm;
  wire mux_190_itm;
  wire mux_209_itm;
  wire mux_232_itm;
  wire mux_246_itm;
  wire mux_272_itm;
  wire mux_340_itm;
  wire mux_351_itm;
  wire mux_378_itm;
  reg weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  reg [7:0] weight_port_read_out_data_0_7_sva;
  reg [7:0] weight_port_read_out_data_0_5_sva;
  reg [14:0] pe_manager_base_bias_sva;
  reg pe_config_is_cluster_sva;
  reg pe_config_is_bias_sva;
  reg [3:0] pe_config_manager_counter_sva;
  reg [7:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8;
  reg [127:0] input_mem_banks_bank_a_0_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_1_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_2_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_3_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_4_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_5_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_6_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_7_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_8_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_9_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_10_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_11_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_12_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_13_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_14_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_15_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_16_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_17_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_18_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_19_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_20_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_21_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_22_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_23_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_24_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_25_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_26_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_27_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_28_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_29_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_30_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_31_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_32_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_33_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_34_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_35_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_36_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_37_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_38_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_39_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_40_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_41_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_42_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_43_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_44_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_45_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_46_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_47_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_48_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_49_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_50_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_51_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_52_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_53_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_54_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_55_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_56_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_57_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_58_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_59_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_60_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_61_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_62_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_63_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_64_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_65_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_66_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_67_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_68_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_69_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_70_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_71_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_72_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_73_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_74_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_75_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_76_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_77_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_78_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_79_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_80_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_81_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_82_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_83_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_84_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_85_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_86_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_87_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_88_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_89_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_90_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_91_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_92_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_93_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_94_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_95_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_96_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_97_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_98_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_99_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_100_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_101_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_102_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_103_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_104_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_105_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_106_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_107_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_108_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_109_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_110_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_111_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_112_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_113_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_114_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_115_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_116_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_117_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_118_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_119_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_120_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_121_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_122_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_123_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_124_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_125_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_126_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_127_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_128_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_129_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_130_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_131_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_132_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_133_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_134_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_135_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_136_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_137_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_138_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_139_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_140_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_141_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_142_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_143_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_144_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_145_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_146_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_147_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_148_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_149_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_150_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_151_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_152_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_153_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_154_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_155_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_156_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_157_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_158_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_159_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_160_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_161_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_162_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_163_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_164_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_165_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_166_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_167_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_168_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_169_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_170_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_171_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_172_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_173_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_174_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_175_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_176_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_177_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_178_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_179_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_180_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_181_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_182_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_183_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_184_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_185_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_186_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_187_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_188_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_189_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_190_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_191_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_192_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_193_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_194_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_195_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_196_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_197_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_198_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_199_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_200_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_201_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_202_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_203_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_204_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_205_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_206_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_207_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_208_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_209_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_210_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_211_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_212_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_213_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_214_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_215_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_216_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_217_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_218_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_219_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_220_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_221_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_222_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_223_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_224_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_225_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_226_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_227_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_228_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_229_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_230_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_231_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_232_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_233_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_234_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_235_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_236_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_237_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_238_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_239_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_240_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_241_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_242_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_243_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_244_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_245_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_246_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_247_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_248_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_249_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_250_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_251_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_252_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_253_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_254_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_255_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_0_6_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_0_8_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_0_9_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_0_11_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_0_12_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_1_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_8_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_9_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_10_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_11_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_12_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_13_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_15_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_8_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_9_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_10_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_11_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_12_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_13_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_4_15_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_8_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_9_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_10_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_11_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_12_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_13_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_14_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_5_15_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_6_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_8_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_9_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_10_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_11_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_12_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_13_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_15_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_0_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_1_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_2_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_3_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_4_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_5_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_6_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_7_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_8_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_9_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_10_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_11_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_12_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_13_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_14_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_15_sva_dfm_1_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_6;
  reg rva_out_reg_data_24_sva_dfm_6;
  reg rva_out_reg_data_31_sva_dfm_6;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_6;
  reg rva_out_reg_data_16_sva_dfm_6;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_6;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_6;
  reg rva_out_reg_data_8_sva_dfm_6;
  reg rva_out_reg_data_0_sva_dfm_6;
  reg [127:0] weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_6;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_6;
  reg [7:0] rva_out_reg_data_103_96_sva_dfm_6;
  reg [7:0] rva_out_reg_data_95_88_sva_dfm_6;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_6;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_6;
  reg rva_out_reg_data_63_sva_dfm_6;
  reg [30:0] accum_vector_data_7_sva_4;
  reg [30:0] accum_vector_data_7_sva_5;
  reg [30:0] accum_vector_data_7_sva_6;
  reg [30:0] accum_vector_data_7_sva_7;
  reg [30:0] accum_vector_data_7_sva_8;
  reg [30:0] accum_vector_data_7_sva_9;
  reg [30:0] accum_vector_data_6_sva_4;
  reg [30:0] accum_vector_data_6_sva_5;
  reg [30:0] accum_vector_data_6_sva_6;
  reg [30:0] accum_vector_data_6_sva_7;
  reg [30:0] accum_vector_data_6_sva_8;
  reg [30:0] accum_vector_data_6_sva_9;
  reg [30:0] accum_vector_data_5_sva_4;
  reg [30:0] accum_vector_data_5_sva_5;
  reg [30:0] accum_vector_data_5_sva_6;
  reg [30:0] accum_vector_data_5_sva_7;
  reg [30:0] accum_vector_data_5_sva_8;
  reg [30:0] accum_vector_data_5_sva_9;
  reg [30:0] accum_vector_data_4_sva_4;
  reg [30:0] accum_vector_data_4_sva_5;
  reg [30:0] accum_vector_data_4_sva_6;
  reg [30:0] accum_vector_data_4_sva_7;
  reg [30:0] accum_vector_data_4_sva_8;
  reg [30:0] accum_vector_data_4_sva_9;
  reg [30:0] accum_vector_data_3_sva_4;
  reg [30:0] accum_vector_data_3_sva_5;
  reg [30:0] accum_vector_data_3_sva_6;
  reg [30:0] accum_vector_data_3_sva_7;
  reg [30:0] accum_vector_data_3_sva_8;
  reg [30:0] accum_vector_data_3_sva_9;
  reg [30:0] accum_vector_data_2_sva_4;
  reg [30:0] accum_vector_data_2_sva_5;
  reg [30:0] accum_vector_data_2_sva_6;
  reg [30:0] accum_vector_data_2_sva_7;
  reg [30:0] accum_vector_data_2_sva_8;
  reg [30:0] accum_vector_data_2_sva_9;
  reg [30:0] accum_vector_data_1_sva_4;
  reg [30:0] accum_vector_data_1_sva_5;
  reg [30:0] accum_vector_data_1_sva_6;
  reg [30:0] accum_vector_data_1_sva_7;
  reg [30:0] accum_vector_data_1_sva_8;
  reg [30:0] accum_vector_data_1_sva_9;
  reg [30:0] accum_vector_data_0_sva_4;
  reg [30:0] accum_vector_data_0_sva_5;
  reg [30:0] accum_vector_data_0_sva_6;
  reg [30:0] accum_vector_data_0_sva_7;
  reg [30:0] accum_vector_data_0_sva_8;
  reg [30:0] accum_vector_data_0_sva_9;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2;
  reg [3:0] pe_config_manager_counter_sva_dfm_3_1;
  reg [7:0] input_read_addrs_sva_1_1;
  wire [8:0] nl_input_read_addrs_sva_1_1;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4_2;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4_3;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4_2;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4_3;
  reg [7:0] rva_out_reg_data_95_88_sva_dfm_4_2;
  reg [7:0] rva_out_reg_data_95_88_sva_dfm_4_3;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4_1;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4_2;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4_3;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_2;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_3;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_1;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_2;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_3;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_3;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_1;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_2;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_4;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_7;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_8;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_9;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_1;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_2;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_5;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_6;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_7;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_2;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_5;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_6_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_7;
  reg [7:0] pe_config_output_counter_sva_dfm_1;
  reg [7:0] pe_config_input_counter_sva_dfm_1;
  reg [127:0] rva_in_reg_data_sva_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_8_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_9_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_10_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_11_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_12_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_13_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_14_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_15_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_2;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_1;
  reg [127:0] input_mem_banks_read_read_data_lpi_1_dfm_1_2;
  reg [127:0] input_mem_banks_read_read_data_lpi_1_dfm_1_3;
  reg [10:0] PEManager_15U_GetWeightAddr_else_acc_3_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_2;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_5;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_6;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_7;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_9;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  reg [14:0] pe_manager_base_weight_sva_dfm_3_1;
  reg [14:0] pe_manager_base_input_sva_dfm_3_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_15_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4;
  reg [7:0] weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1;
  reg [7:0] weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_14_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_30_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_30_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_44_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_1;
  reg weight_mem_run_3_for_5_and_148_itm_1;
  reg weight_mem_run_3_for_5_and_148_itm_2;
  reg weight_mem_run_3_for_5_and_150_itm_1;
  reg weight_mem_run_3_for_5_and_150_itm_2;
  reg weight_mem_run_3_for_5_and_7_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
  reg weight_mem_run_3_for_5_and_12_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_2;
  reg weight_mem_run_3_for_5_and_28_itm_1;
  reg weight_mem_run_3_for_5_and_28_itm_2;
  reg weight_mem_run_3_for_5_and_30_itm_1;
  reg weight_mem_run_3_for_5_and_30_itm_2;
  reg weight_mem_run_3_for_5_and_31_itm_1;
  reg weight_mem_run_3_for_5_and_31_itm_2;
  reg weight_mem_run_3_for_5_and_100_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1;
  reg weight_mem_run_3_for_5_and_135_itm_1;
  reg weight_mem_run_3_for_5_and_136_itm_1;
  reg weight_mem_run_3_for_5_and_142_itm_1;
  reg ProductSum_for_asn_128_itm_2;
  reg ProductSum_for_asn_128_itm_4;
  reg ProductSum_for_asn_108_itm_2;
  reg ProductSum_for_asn_108_itm_4;
  reg ProductSum_for_asn_95_itm_1;
  reg ProductSum_for_asn_95_itm_2;
  reg ProductSum_for_asn_95_itm_3;
  reg ProductSum_for_asn_95_itm_4;
  reg ProductSum_for_asn_95_itm_5;
  reg ProductSum_for_asn_82_itm_1;
  reg ProductSum_for_asn_82_itm_2;
  reg ProductSum_for_asn_82_itm_3;
  reg ProductSum_for_asn_82_itm_4;
  reg ProductSum_for_asn_69_itm_1;
  reg ProductSum_for_asn_69_itm_2;
  reg ProductSum_for_asn_69_itm_4;
  reg ProductSum_for_asn_69_itm_5;
  reg ProductSum_for_asn_56_itm_2;
  reg ProductSum_for_asn_56_itm_4;
  reg ProductSum_for_asn_41_itm_2;
  reg ProductSum_for_asn_41_itm_4;
  reg ProductSum_for_asn_28_itm_2;
  reg ProductSum_for_asn_28_itm_4;
  reg accum_vector_operator_1_for_asn_10_itm_7;
  reg accum_vector_operator_1_for_asn_13_itm_2;
  reg accum_vector_operator_1_for_asn_13_itm_3;
  reg accum_vector_operator_1_for_asn_13_itm_4;
  reg accum_vector_operator_1_for_asn_13_itm_5;
  reg accum_vector_operator_1_for_asn_13_itm_6;
  reg accum_vector_operator_1_for_asn_25_itm_7;
  reg accum_vector_operator_1_for_asn_28_itm_3;
  reg accum_vector_operator_1_for_asn_28_itm_4;
  reg accum_vector_operator_1_for_asn_28_itm_5;
  reg accum_vector_operator_1_for_asn_28_itm_6;
  reg accum_vector_operator_1_for_asn_43_itm_3;
  reg accum_vector_operator_1_for_asn_43_itm_4;
  reg accum_vector_operator_1_for_asn_43_itm_5;
  reg accum_vector_operator_1_for_asn_43_itm_6;
  reg accum_vector_operator_1_for_asn_43_itm_7;
  reg accum_vector_operator_1_for_asn_55_itm_7;
  reg accum_vector_operator_1_for_asn_58_itm_2;
  reg accum_vector_operator_1_for_asn_58_itm_3;
  reg accum_vector_operator_1_for_asn_58_itm_4;
  reg accum_vector_operator_1_for_asn_58_itm_5;
  reg accum_vector_operator_1_for_asn_58_itm_6;
  reg accum_vector_operator_1_for_asn_73_itm_3;
  reg accum_vector_operator_1_for_asn_73_itm_4;
  reg accum_vector_operator_1_for_asn_73_itm_5;
  reg accum_vector_operator_1_for_asn_73_itm_6;
  reg accum_vector_operator_1_for_asn_73_itm_7;
  reg accum_vector_operator_1_for_asn_85_itm_7;
  reg accum_vector_operator_1_for_asn_88_itm_1;
  reg accum_vector_operator_1_for_asn_88_itm_2;
  reg accum_vector_operator_1_for_asn_88_itm_3;
  reg accum_vector_operator_1_for_asn_88_itm_4;
  reg accum_vector_operator_1_for_asn_88_itm_5;
  reg accum_vector_operator_1_for_asn_88_itm_6;
  reg accum_vector_operator_1_for_asn_100_itm_7;
  reg accum_vector_operator_1_for_asn_103_itm_2;
  reg accum_vector_operator_1_for_asn_103_itm_3;
  reg accum_vector_operator_1_for_asn_103_itm_4;
  reg accum_vector_operator_1_for_asn_103_itm_5;
  reg accum_vector_operator_1_for_asn_103_itm_6;
  reg accum_vector_operator_1_for_asn_115_itm_7;
  reg accum_vector_operator_1_for_asn_118_itm_2;
  reg accum_vector_operator_1_for_asn_118_itm_3;
  reg accum_vector_operator_1_for_asn_118_itm_4;
  reg accum_vector_operator_1_for_asn_118_itm_5;
  reg accum_vector_operator_1_for_asn_118_itm_6;
  reg [14:0] PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1;
  reg while_if_mux_27_itm_1;
  reg PECore_PushAxiRsp_mux_10_itm_1;
  reg PECore_PushAxiRsp_mux_23_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
  reg [119:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_8;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_3_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0;
  wire [30:0] accum_vector_data_7_sva_8_mx0w0;
  wire [30:0] accum_vector_data_7_sva_7_mx0w0;
  wire [30:0] accum_vector_data_7_sva_6_mx0w0;
  wire [30:0] accum_vector_data_7_sva_5_mx0w0;
  wire [30:0] accum_vector_data_7_sva_4_mx0w0;
  wire [30:0] accum_vector_data_6_sva_8_mx0w0;
  wire [30:0] accum_vector_data_6_sva_7_mx0w0;
  wire [30:0] accum_vector_data_6_sva_6_mx0w0;
  wire [30:0] accum_vector_data_6_sva_5_mx0w0;
  wire [30:0] accum_vector_data_6_sva_4_mx0w0;
  wire [30:0] accum_vector_data_5_sva_8_mx0w0;
  wire [30:0] accum_vector_data_5_sva_7_mx0w0;
  wire [30:0] accum_vector_data_5_sva_6_mx0w0;
  wire [30:0] accum_vector_data_5_sva_5_mx0w0;
  wire [30:0] accum_vector_data_5_sva_4_mx0w0;
  wire [30:0] accum_vector_data_4_sva_9_mx0w0;
  wire [30:0] accum_vector_data_4_sva_8_mx0w0;
  wire [30:0] accum_vector_data_4_sva_7_mx0w0;
  wire [30:0] accum_vector_data_4_sva_6_mx0w0;
  wire [30:0] accum_vector_data_4_sva_5_mx0w0;
  wire [30:0] accum_vector_data_4_sva_4_mx0w0;
  wire [30:0] accum_vector_data_3_sva_8_mx0w0;
  wire [30:0] accum_vector_data_3_sva_7_mx0w0;
  wire [30:0] accum_vector_data_3_sva_6_mx0w0;
  wire [30:0] accum_vector_data_3_sva_5_mx0w0;
  wire [30:0] accum_vector_data_3_sva_4_mx0w0;
  wire [30:0] accum_vector_data_2_sva_9_mx0w0;
  wire [30:0] accum_vector_data_2_sva_8_mx0w0;
  wire [30:0] accum_vector_data_2_sva_7_mx0w0;
  wire [30:0] accum_vector_data_2_sva_6_mx0w0;
  wire [30:0] accum_vector_data_2_sva_5_mx0w0;
  wire [30:0] accum_vector_data_2_sva_4_mx0w0;
  wire [30:0] accum_vector_data_1_sva_8_mx0w0;
  wire [30:0] accum_vector_data_1_sva_7_mx0w0;
  wire [30:0] accum_vector_data_1_sva_6_mx0w0;
  wire [30:0] accum_vector_data_1_sva_5_mx0w0;
  wire [30:0] accum_vector_data_1_sva_4_mx0w0;
  wire [30:0] accum_vector_data_0_sva_8_mx0w0;
  wire [30:0] accum_vector_data_0_sva_7_mx0w0;
  wire [30:0] accum_vector_data_0_sva_6_mx0w0;
  wire [30:0] accum_vector_data_0_sva_5_mx0w0;
  wire [30:0] accum_vector_data_0_sva_4_mx0w0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_39_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_38_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_37_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0;
  wire weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_12_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_11_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_8_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_4_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_3_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0;
  wire [14:0] weight_read_addrs_1_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_3_lpi_1_dfm_1_1;
  wire [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_5_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_7_lpi_1_dfm_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  wire accum_vector_data_3_sva_1_load_mx0w1;
  wire [7:0] pe_config_output_counter_sva_mx1;
  wire pe_config_is_zero_first_sva_mx1;
  wire pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  wire [7:0] weight_port_read_out_data_0_7_sva_mx0;
  wire [7:0] weight_port_read_out_data_0_5_sva_mx0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
  wire [7:0] weight_port_read_out_data_0_7_sva_dfm_mx0w1;
  wire [7:0] weight_port_read_out_data_0_5_sva_dfm_mx0w1;
  wire PECore_PushAxiRsp_if_else_mux_10_mx0w2;
  wire PECore_PushAxiRsp_if_else_mux_23_mx0w2;
  wire [7:0] rva_out_reg_data_103_96_sva_dfm_4_mx0w0;
  wire [7:0] rva_out_reg_data_95_88_sva_dfm_4_mx0w0;
  wire [7:0] rva_out_reg_data_79_72_sva_dfm_4_mx0w0;
  wire [7:0] rva_out_reg_data_71_64_sva_dfm_4_mx0w0;
  wire rva_out_reg_data_63_sva_dfm_6_mx1;
  wire [7:0] rva_out_reg_data_55_48_sva_dfm_6_mx1;
  wire [6:0] rva_out_reg_data_62_56_sva_dfm_6_mx1;
  wire [6:0] rva_out_reg_data_46_40_sva_dfm_6_mx1;
  wire [3:0] rva_out_reg_data_39_36_sva_dfm_6_mx1;
  wire [3:0] rva_out_reg_data_35_32_sva_dfm_6_mx1;
  wire accum_vector_data_5_sva_1_load_mx0w0;
  wire input_read_req_valid_lpi_1_dfm_1_mx0w2;
  wire [14:0] pe_manager_base_input_sva_mx2;
  wire accum_vector_data_7_sva_1_load_mx0w1;
  wire accum_vector_data_6_sva_1_load_mx0w1;
  wire accum_vector_data_1_sva_1_load_mx0w1;
  wire accum_vector_data_0_sva_1_load_mx0w1;
  wire accum_vector_data_4_sva_1_load_mx0w0;
  wire accum_vector_data_2_sva_1_load_mx0w0;
  wire PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_4;
  wire while_and_1266_cse_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
  wire [7:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1;
  wire weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_sva_1;
  wire rva_out_reg_data_63_sva_dfm_7;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
  wire PECore_PushAxiRsp_if_asn_79;
  wire PECore_PushAxiRsp_if_asn_81;
  wire PECore_PushAxiRsp_if_asn_83;
  wire weight_mem_run_3_for_5_asn_447;
  wire weight_mem_run_3_for_5_asn_449;
  wire weight_mem_run_3_for_5_asn_451;
  wire weight_mem_run_3_for_5_asn_453;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434;
  wire PECore_PushAxiRsp_if_asn_87;
  wire PECore_PushAxiRsp_if_asn_89;
  wire PECore_PushAxiRsp_if_asn_91;
  wire while_asn_998;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367;
  wire weight_mem_run_3_for_5_and_152;
  wire weight_mem_run_3_for_5_and_156;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371;
  wire [7:0] pe_manager_base_input_sva_mx1_7_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0;
  wire mux_136_cse;
  wire PECore_PushAxiRsp_if_mux1h_15;
  wire [5:0] PECore_PushAxiRsp_if_mux1h_16;
  wire PECore_PushAxiRsp_if_mux1h_17;
  wire [7:0] weight_port_read_out_data_7_0_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_3_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_2_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_5_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_4_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_7_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_6_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_9_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_8_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_11_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_10_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_13_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_12_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_15_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_7_14_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_5_15_sva_dfm_1_2;
  wire [7:0] weight_port_read_out_data_5_14_sva_dfm_1_2;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse;
  reg reg_rva_in_reg_rw_sva_2_cse;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2;
  reg reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse;
  wire nor_329_cse;
  reg [1:0] weight_mem_run_3_for_5_mux_109_itm_1_7_6;
  reg [5:0] weight_mem_run_3_for_5_mux_109_itm_1_5_0;
  wire weight_mem_run_3_for_5_and_199_ssc;
  reg weight_mem_run_3_for_5_mux_107_itm_1_7;
  reg [6:0] weight_mem_run_3_for_5_mux_107_itm_1_6_0;
  reg weight_mem_run_3_for_5_mux_110_itm_1_7;
  reg [6:0] weight_mem_run_3_for_5_mux_110_itm_1_6_0;
  wire weight_mem_run_3_for_5_and_202_ssc;
  reg weight_mem_run_3_for_5_mux_111_itm_1_7;
  reg [6:0] weight_mem_run_3_for_5_mux_111_itm_1_6_0;
  reg weight_mem_run_3_for_5_mux_108_itm_1_7;
  reg [6:0] weight_mem_run_3_for_5_mux_108_itm_1_6_0;
  reg weight_mem_run_3_for_5_mux_11_itm_1_7;
  reg [6:0] weight_mem_run_3_for_5_mux_11_itm_1_6_0;
  reg [1:0] weight_mem_run_3_for_5_mux_12_itm_1_7_6;
  reg [5:0] weight_mem_run_3_for_5_mux_12_itm_1_5_0;
  wire weight_mem_banks_load_store_for_else_and_ssc;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_7_4;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_3_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0;
  wire weight_mem_banks_load_store_for_else_and_3_ssc;
  reg [1:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7_6;
  reg [5:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_5_0;
  wire weight_mem_banks_load_store_for_else_and_77_ssc;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7_4;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_3_0;
  reg weight_port_read_out_data_0_3_sva_dfm_1_7;
  reg [6:0] weight_port_read_out_data_0_3_sva_dfm_1_6_0;
  wire and_1022_ssc;
  reg weight_port_read_out_data_0_2_sva_dfm_1_7;
  reg [6:0] weight_port_read_out_data_0_2_sva_dfm_1_6_0;
  wire weight_port_read_out_data_and_136_ssc;
  reg [3:0] weight_port_read_out_data_0_1_sva_dfm_1_7_4;
  reg [3:0] weight_port_read_out_data_0_1_sva_dfm_1_3_0;
  wire and_1042_ssc;
  wire [3:0] weight_port_read_out_data_0_0_sva_dfm_mx0w1_7_4;
  wire [3:0] weight_port_read_out_data_0_0_sva_dfm_mx0w1_3_0;
  wire [1:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000;
  wire [5:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000001;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000;
  wire [6:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000;
  wire [6:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001;
  reg [3:0] weight_port_read_out_data_0_1_sva_dfm_2_rsp_0;
  reg [3:0] weight_port_read_out_data_0_1_sva_dfm_2_rsp_1;
  reg weight_port_read_out_data_0_2_sva_dfm_2_rsp_0;
  reg [6:0] weight_port_read_out_data_0_2_sva_dfm_2_rsp_1;
  reg weight_port_read_out_data_0_3_sva_dfm_2_rsp_0;
  reg [6:0] weight_port_read_out_data_0_3_sva_dfm_2_rsp_1;
  reg [3:0] reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd;
  reg [3:0] reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd;
  reg [6:0] reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_1;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd;
  reg [6:0] reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd_1;
  wire [3:0] weight_port_read_out_data_0_1_sva_mx0_7_4;
  wire [3:0] weight_port_read_out_data_0_1_sva_mx0_3_0;
  wire weight_port_read_out_data_and_129_ssc;
  reg [3:0] weight_port_read_out_data_0_0_sva_dfm_1_1_7_4;
  reg [3:0] weight_port_read_out_data_0_0_sva_dfm_1_1_3_0;
  wire weight_port_read_out_data_0_3_sva_mx0_7;
  wire [6:0] weight_port_read_out_data_0_3_sva_mx0_6_0;
  wire weight_port_read_out_data_0_2_sva_mx0_7;
  wire [6:0] weight_port_read_out_data_0_2_sva_mx0_6_0;
  reg [3:0] weight_port_read_out_data_0_0_sva_dfm_2_7_4;
  reg [3:0] weight_port_read_out_data_0_0_sva_dfm_2_3_0;
  reg weight_port_read_out_data_0_13_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_13_sva_dfm_2_6_0;
  reg weight_port_read_out_data_0_14_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_14_sva_dfm_2_6_0;
  reg [1:0] weight_port_read_out_data_0_15_sva_dfm_2_7_6;
  reg [5:0] weight_port_read_out_data_0_15_sva_dfm_2_5_0;
  wire [1:0] rva_out_reg_data_127_120_sva_dfm_4_mx0w0_7_6;
  wire [5:0] rva_out_reg_data_127_120_sva_dfm_4_mx0w0_5_0;
  wire rva_out_reg_data_119_112_sva_dfm_4_mx0w0_7;
  wire [6:0] rva_out_reg_data_119_112_sva_dfm_4_mx0w0_6_0;
  wire rva_out_reg_data_111_104_sva_dfm_4_mx0w0_7;
  wire [6:0] rva_out_reg_data_111_104_sva_dfm_4_mx0w0_6_0;
  reg rva_out_reg_data_111_104_sva_dfm_4_1_7;
  reg [6:0] rva_out_reg_data_111_104_sva_dfm_4_1_6_0;
  reg rva_out_reg_data_119_112_sva_dfm_4_1_7;
  reg [6:0] rva_out_reg_data_119_112_sva_dfm_4_1_6_0;
  wire rva_out_reg_data_and_78_ssc;
  reg [1:0] rva_out_reg_data_127_120_sva_dfm_4_1_7_6;
  reg [5:0] rva_out_reg_data_127_120_sva_dfm_4_1_5_0;
  wire weight_mem_run_3_for_5_and_165_ssc;
  wire weight_mem_run_3_for_5_and_166_ssc;
  wire weight_mem_run_3_for_5_and_168_ssc;
  wire weight_mem_run_3_for_5_and_170_ssc;
  wire weight_mem_run_3_for_5_and_171_ssc;
  reg weight_port_read_out_data_0_2_sva_dfm_1_1_7;
  reg [6:0] weight_port_read_out_data_0_2_sva_dfm_1_1_6_0;
  wire weight_mem_run_3_for_5_and_157_ssc;
  wire weight_mem_run_3_for_5_and_158_ssc;
  wire weight_mem_run_3_for_5_and_160_ssc;
  wire weight_mem_run_3_for_5_and_162_ssc;
  wire weight_mem_run_3_for_5_and_163_ssc;
  wire weight_port_read_out_data_and_130_ssc;
  reg weight_port_read_out_data_0_3_sva_dfm_1_1_7;
  reg [6:0] weight_port_read_out_data_0_3_sva_dfm_1_1_6_0;
  reg weight_mem_run_3_for_5_mux_13_itm_1_7;
  reg [6:0] weight_mem_run_3_for_5_mux_13_itm_1_6_0;
  reg weight_mem_run_3_for_5_mux_14_itm_1_7;
  reg [6:0] weight_mem_run_3_for_5_mux_14_itm_1_6_0;
  reg [1:0] weight_mem_run_3_for_5_mux_15_itm_1_7_6;
  reg [5:0] weight_mem_run_3_for_5_mux_15_itm_1_5_0;
  reg weight_port_read_out_data_0_3_sva_7;
  reg [6:0] weight_port_read_out_data_0_3_sva_6_0;
  reg weight_port_read_out_data_0_2_sva_7;
  reg [6:0] weight_port_read_out_data_0_2_sva_6_0;
  reg [3:0] weight_port_read_out_data_0_1_sva_7_4;
  reg [3:0] weight_port_read_out_data_0_1_sva_3_0;
  reg [1:0] rva_out_reg_data_127_120_sva_dfm_6_7_6;
  reg [5:0] rva_out_reg_data_127_120_sva_dfm_6_5_0;
  reg rva_out_reg_data_119_112_sva_dfm_6_7;
  reg [6:0] rva_out_reg_data_119_112_sva_dfm_6_6_0;
  reg rva_out_reg_data_111_104_sva_dfm_6_7;
  reg [6:0] rva_out_reg_data_111_104_sva_dfm_6_6_0;
  wire and_568_ssc;
  wire and_569_ssc;
  wire and_570_ssc;
  reg [3:0] weight_port_read_out_data_0_1_sva_dfm_1_1_7_4;
  reg [3:0] weight_port_read_out_data_0_1_sva_dfm_1_1_3_0;
  reg weight_port_read_out_data_0_3_sva_dfm_4_7;
  reg [6:0] weight_port_read_out_data_0_3_sva_dfm_4_6_0;
  wire weight_port_read_out_data_and_209_ssc;
  reg [3:0] weight_port_read_out_data_0_0_sva_dfm_2_7_4_1;
  reg [3:0] weight_port_read_out_data_0_0_sva_dfm_2_3_0_1;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_6;
  reg [5:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_5_0;
  reg [3:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_6_3;
  reg [2:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_2_0;
  wire [3:0] weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_7_4;
  wire [3:0] weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_3_0;
  wire rva_out_reg_data_and_23_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_2_cse;
  wire rva_out_reg_data_and_26_cse;
  wire input_mem_banks_read_read_data_and_cse;
  wire weight_port_read_out_data_and_122_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_cse;
  wire PECore_RunScale_if_and_cse;
  wire rva_in_reg_rw_and_cse;
  wire accum_vector_operator_1_for_and_cse;
  wire ProductSum_for_and_cse;
  wire data_in_tmp_operator_2_for_and_cse;
  wire weight_mem_run_3_for_aelse_and_cse;
  wire data_in_tmp_operator_2_for_and_16_cse;
  wire weight_mem_banks_read_1_read_data_and_8_cse;
  wire ProductSum_for_and_8_cse;
  wire weight_mem_run_3_for_aelse_and_4_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_375_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_380_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_382_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_cse;
  wire weight_read_addrs_and_5_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_2_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_4_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_48_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_54_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_60_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_66_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_72_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_78_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_84_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_90_cse;
  wire weight_read_addrs_and_7_cse;
  wire weight_write_data_data_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_15_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_22_cse;
  wire Arbiter_8U_Roundrobin_pick_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_25_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_64_cse;
  wire weight_write_data_data_and_16_cse;
  wire PECore_DecodeAxiWrite_switch_lp_and_2_cse;
  wire rva_in_reg_rw_and_5_cse;
  wire PECore_UpdateFSM_switch_lp_and_9_cse;
  wire state_and_cse;
  wire PECore_PushOutput_if_and_cse;
  wire weight_port_read_out_data_and_138_cse;
  wire PECore_RunMac_if_and_2_cse;
  wire weight_read_addrs_and_17_cse;
  wire weight_port_read_out_data_and_143_cse;
  wire weight_port_read_out_data_and_158_cse;
  wire weight_port_read_out_data_and_137_cse;
  wire weight_port_read_out_data_and_185_cse;
  wire weight_port_read_out_data_and_199_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_384_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_379_cse;
  wire while_if_and_10_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_30_cse;
  wire rva_in_reg_rw_and_2_cse;
  wire ProductSum_for_and_14_cse;
  wire weight_read_addrs_and_19_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_404_cse;
  wire weight_read_addrs_and_20_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_408_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_152_cse;
  wire input_mem_banks_read_read_data_and_9_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse;
  wire while_if_and_14_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_7_cse;
  wire while_if_and_6_cse;
  wire rva_out_reg_data_and_41_cse;
  wire input_read_req_valid_and_1_cse;
  wire weight_mem_banks_load_store_for_else_and_4_cse;
  wire weight_mem_banks_load_store_for_else_and_1_cse;
  wire weight_mem_banks_load_store_for_else_and_2_cse;
  wire weight_mem_banks_load_store_for_else_and_56_cse;
  wire weight_mem_banks_load_store_for_else_and_57_cse;
  wire weight_mem_banks_load_store_for_else_and_62_cse;
  wire weight_mem_banks_load_store_for_else_and_67_cse;
  wire weight_mem_banks_load_store_for_else_and_64_cse;
  wire rva_in_reg_rw_and_6_cse;
  wire rva_in_reg_rw_and_7_cse;
  wire PECore_RunMac_if_and_3_cse;
  wire ProductSum_for_and_22_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_410_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_158_cse;
  wire input_mem_banks_read_read_data_and_18_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse;
  wire ProductSum_for_and_26_cse;
  wire pe_manager_base_weight_and_5_cse;
  wire pe_manager_base_weight_and_6_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_11_cse;
  wire while_if_and_7_cse;
  wire rva_out_reg_data_and_57_cse;
  wire input_read_req_valid_and_2_cse;
  wire weight_mem_read_arbxbar_xbar_requests_transpose_and_13_cse;
  wire rva_in_reg_rw_and_10_cse;
  wire ProductSum_for_and_30_cse;
  wire input_mem_banks_read_read_data_and_27_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_15_cse;
  wire input_read_req_valid_and_3_cse;
  wire rva_out_reg_data_and_93_cse;
  wire rva_in_reg_rw_and_3_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_19_cse;
  wire PECore_RunMac_if_and_10_cse;
  wire accum_vector_operator_1_for_and_45_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_23_cse;
  wire rva_out_reg_data_and_101_cse;
  wire rva_out_reg_data_and_104_cse;
  wire PECore_RunMac_if_and_8_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse;
  wire rva_out_reg_data_and_109_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_29_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_35_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_40_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse;
  wire act_port_reg_data_and_16_cse;
  reg [3:0] weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
  reg [3:0] weight_port_read_out_data_0_0_sva_dfm_3_rsp_1;
  reg [1:0] rva_out_reg_data_127_120_sva_dfm_4_2_rsp_0;
  reg [5:0] rva_out_reg_data_127_120_sva_dfm_4_2_rsp_1;
  reg rva_out_reg_data_119_112_sva_dfm_4_2_rsp_0;
  reg [6:0] rva_out_reg_data_119_112_sva_dfm_4_2_rsp_1;
  reg rva_out_reg_data_111_104_sva_dfm_4_2_rsp_0;
  reg [6:0] rva_out_reg_data_111_104_sva_dfm_4_2_rsp_1;
  reg [3:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd;
  reg [2:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1;
  reg [1:0] reg_rva_out_reg_data_127_120_sva_dfm_4_3_ftd;
  reg [5:0] reg_rva_out_reg_data_127_120_sva_dfm_4_3_ftd_1;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd;
  reg [6:0] reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd_1;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd;
  reg [6:0] reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd_1;
  wire [3:0] weight_port_read_out_data_0_4_sva_mx0_7_4;
  wire [3:0] weight_port_read_out_data_0_4_sva_mx0_3_0;
  wire [3:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000000;
  wire [3:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000001;
  wire rva_out_reg_data_111_104_sva_dfm_7_7;
  wire rva_out_reg_data_119_112_sva_dfm_7_7;
  wire [1:0] rva_out_reg_data_127_120_sva_dfm_7_7_6;
  wire [3:0] PECore_PushAxiRsp_if_mux1h_12_6_3;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_12_2_0;
  wire PECore_PushAxiRsp_if_mux1h_14_6;
  wire [5:0] PECore_PushAxiRsp_if_mux1h_14_5_0;
  reg [1:0] rva_out_reg_data_127_120_sva_dfm_4_4_7_6;
  reg [5:0] rva_out_reg_data_127_120_sva_dfm_4_4_5_0;
  reg rva_out_reg_data_119_112_sva_dfm_4_4_7;
  reg [6:0] rva_out_reg_data_119_112_sva_dfm_4_4_6_0;
  reg rva_out_reg_data_111_104_sva_dfm_4_4_7;
  reg [6:0] rva_out_reg_data_111_104_sva_dfm_4_4_6_0;
  wire weight_mem_run_3_for_5_and_187_ssc;
  reg [3:0] weight_port_read_out_data_0_4_sva_dfm_1_1_7_4;
  reg [3:0] weight_port_read_out_data_0_4_sva_dfm_1_1_3_0;
  reg [3:0] weight_port_read_out_data_0_4_sva_7_4;
  reg [3:0] weight_port_read_out_data_0_4_sva_3_0;
  reg [3:0] weight_port_read_out_data_0_10_sva_dfm_2_7_4;
  reg [3:0] weight_port_read_out_data_0_10_sva_dfm_2_3_0;
  reg rva_out_reg_data_23_17_sva_dfm_6_6;
  reg [5:0] rva_out_reg_data_23_17_sva_dfm_6_5_0;
  reg [3:0] rva_out_reg_data_15_9_sva_dfm_6_6_3;
  reg [2:0] rva_out_reg_data_15_9_sva_dfm_6_2_0;
  wire and_1050_ssc;
  wire and_1052_ssc;
  wire and_1053_ssc;
  wire [3:0] weight_port_read_out_data_0_4_sva_dfm_mx0w2_7_4;
  wire [3:0] weight_port_read_out_data_0_4_sva_dfm_mx0w2_3_0;
  wire [3:0] rva_out_reg_data_87_80_sva_dfm_4_mx0w0_7_4;
  wire [3:0] rva_out_reg_data_87_80_sva_dfm_4_mx0w0_3_0;
  wire [3:0] PECore_PushAxiRsp_if_mux1h_10_6_3;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_10_2_0;
  reg [3:0] rva_out_reg_data_7_1_sva_dfm_6_rsp_0;
  reg [2:0] rva_out_reg_data_7_1_sva_dfm_6_rsp_1;
  reg [3:0] rva_out_reg_data_87_80_sva_dfm_4_1_7_4;
  reg [3:0] rva_out_reg_data_87_80_sva_dfm_4_1_3_0;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_1_7_4;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_1_3_0;
  reg [3:0] rva_out_reg_data_87_80_sva_dfm_6_7_4;
  reg [3:0] rva_out_reg_data_87_80_sva_dfm_6_3_0;
  reg [3:0] rva_out_reg_data_87_80_sva_dfm_4_2_7_4;
  reg [3:0] rva_out_reg_data_87_80_sva_dfm_4_2_3_0;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_2_7_4;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_2_3_0;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_3_rsp_0;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_3_rsp_1;
  reg [3:0] rva_out_reg_data_87_80_sva_dfm_4_3_rsp_0;
  reg [3:0] rva_out_reg_data_87_80_sva_dfm_4_3_rsp_1;
  reg [3:0] reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd;
  reg [3:0] reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd_1;
  reg [3:0] reg_rva_out_reg_data_87_80_sva_dfm_4_4_ftd;
  reg [3:0] reg_rva_out_reg_data_87_80_sva_dfm_4_4_ftd_1;
  wire or_tmp_484;
  wire not_tmp_488;
  wire mux_tmp_427;
  wire mux_tmp_429;
  wire and_dcpl_949;
  wire and_dcpl_958;
  wire or_dcpl_390;
  wire or_dcpl_394;
  wire or_dcpl_395;
  wire or_dcpl_403;
  wire or_dcpl_407;
  wire or_dcpl_408;
  wire or_tmp_541;
  wire and_tmp_17;
  wire and_tmp_18;
  wire or_tmp_583;
  wire or_tmp_584;
  wire or_tmp_607;
  wire or_tmp_608;
  wire mux_tmp_512;
  wire mux_tmp_514;
  wire mux_tmp_519;
  wire mux_tmp_548;
  wire and_1125_cse;
  wire and_1140_cse;
  wire and_1155_cse;
  wire and_1170_cse;
  wire and_1188_cse;
  wire and_1203_cse;
  wire and_1221_cse;
  wire and_1236_cse;
  wire or_931_cse;
  wire or_928_cse;
  wire or_945_cse;
  wire nor_571_cse;
  wire and_1279_cse;
  wire xor_1_cse;
  wire and_1327_cse;
  wire mux_468_cse;
  wire and_1397_cse;
  wire and_1442_cse;
  wire and_1463_cse;
  wire or_1098_cse;
  wire or_1097_cse;
  wire nor_589_cse;
  wire and_1287_cse;
  wire and_1600_cse;
  wire nor_573_cse;
  wire nor_582_cse;
  wire nand_91_cse;
  wire nor_524_cse;
  wire nand_76_cse;
  wire and_1607_cse;
  wire and_1608_cse;
  wire and_1332_cse;
  wire and_1352_cse;
  wire and_1488_cse;
  wire and_1557_cse;
  wire act_port_reg_data_act_port_reg_data_nor_cse;
  wire mux_494_cse;
  wire and_1086_cse;
  wire or_939_cse;
  wire and_1363_cse;
  wire mux_87_cse;
  wire and_1551_cse;
  wire and_1580_cse;
  wire mux_522_cse;
  wire and_1529_cse;
  reg reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_79_72_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_71_64_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  reg reg_weight_read_addrs_3_lpi_1_dfm_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2_enexo;
  reg reg_weight_read_addrs_3_lpi_1_dfm_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_enexo_1;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2;
  reg reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2_enexo_1;
  reg reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  reg reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_manager_base_input_enexo;
  reg reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_config_num_output_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_2_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_2_1_enexo;
  reg reg_rva_in_reg_data_sva_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_2_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_127_120_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_79_72_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_71_64_sva_dfm_4_2_enexo;
  reg reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_11_itm_1_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_107_itm_1_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_108_itm_1_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_109_itm_1_1_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_12_itm_1_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_111_itm_1_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_110_itm_1_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_79_72_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_71_64_sva_dfm_4_1_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1;
  reg reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo;
  reg reg_pe_config_input_counter_sva_dfm_1_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_1_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_1_1_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_1_1_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_3_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_3_1_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_3_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_2_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_1_1_1_enexo;
  reg reg_rva_out_reg_data_127_120_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_127_120_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_1_1_enexo;
  wire rva_out_reg_data_and_128_enex5;
  wire rva_out_reg_data_and_129_enex5;
  wire rva_out_reg_data_and_130_enex5;
  wire rva_out_reg_data_and_131_enex5;
  wire rva_out_reg_data_and_132_enex5;
  wire rva_out_reg_data_and_133_enex5;
  wire rva_out_reg_data_and_134_enex5;
  wire rva_out_reg_data_and_135_enex5;
  wire rva_out_reg_data_and_136_enex5;
  wire rva_out_reg_data_and_137_enex5;
  wire rva_out_reg_data_and_138_enex5;
  wire rva_out_reg_data_and_139_enex5;
  wire rva_out_reg_data_and_140_enex5;
  wire rva_out_reg_data_and_141_enex5;
  wire rva_out_reg_data_and_142_enex5;
  wire input_mem_banks_read_read_data_and_35_enex5;
  wire weight_port_read_out_data_and_213_enex5;
  wire input_mem_banks_read_read_data_and_36_enex5;
  wire input_mem_banks_read_read_data_and_37_enex5;
  wire input_mem_banks_read_read_data_and_38_enex5;
  wire input_mem_banks_read_1_read_data_and_enex5;
  wire weight_port_read_out_data_and_214_enex5;
  wire weight_port_read_out_data_and_215_enex5;
  wire weight_port_read_out_data_and_216_enex5;
  wire weight_port_read_out_data_and_217_enex5;
  wire weight_port_read_out_data_and_218_enex5;
  wire weight_port_read_out_data_and_219_enex5;
  wire weight_port_read_out_data_and_220_enex5;
  wire weight_port_read_out_data_and_221_enex5;
  wire weight_port_read_out_data_and_222_enex5;
  wire weight_port_read_out_data_and_223_enex5;
  wire weight_port_read_out_data_and_224_enex5;
  wire weight_port_read_out_data_and_225_enex5;
  wire weight_port_read_out_data_and_226_enex5;
  wire weight_port_read_out_data_and_227_enex5;
  wire weight_port_read_out_data_and_228_enex5;
  wire weight_port_read_out_data_and_15_enex5;
  wire weight_port_read_out_data_and_229_enex5;
  wire weight_port_read_out_data_and_230_enex5;
  wire weight_port_read_out_data_and_231_enex5;
  wire weight_port_read_out_data_and_232_enex5;
  wire weight_port_read_out_data_and_233_enex5;
  wire weight_port_read_out_data_and_234_enex5;
  wire weight_port_read_out_data_and_235_enex5;
  wire weight_port_read_out_data_and_236_enex5;
  wire weight_port_read_out_data_and_237_enex5;
  wire weight_port_read_out_data_and_238_enex5;
  wire weight_port_read_out_data_and_239_enex5;
  wire weight_port_read_out_data_and_240_enex5;
  wire weight_port_read_out_data_and_241_enex5;
  wire weight_port_read_out_data_and_242_enex5;
  wire weight_port_read_out_data_and_243_enex5;
  wire weight_port_read_out_data_and_31_enex5;
  wire input_mem_banks_read_1_read_data_and_5_enex5;
  wire weight_read_addrs_and_28_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5;
  wire weight_write_data_data_and_48_enex5;
  wire weight_write_data_data_and_49_enex5;
  wire weight_write_data_data_and_50_enex5;
  wire weight_write_data_data_and_51_enex5;
  wire weight_write_data_data_and_52_enex5;
  wire weight_write_data_data_and_53_enex5;
  wire weight_write_data_data_and_54_enex5;
  wire weight_write_data_data_and_55_enex5;
  wire weight_write_data_data_and_56_enex5;
  wire weight_write_data_data_and_57_enex5;
  wire weight_write_data_data_and_58_enex5;
  wire weight_write_data_data_and_59_enex5;
  wire weight_write_data_data_and_60_enex5;
  wire weight_write_data_data_and_61_enex5;
  wire weight_write_data_data_and_62_enex5;
  wire weight_write_data_data_and_63_enex5;
  wire weight_write_addrs_and_enex5;
  wire weight_write_data_data_and_64_enex5;
  wire weight_write_data_data_and_65_enex5;
  wire weight_write_data_data_and_66_enex5;
  wire weight_write_data_data_and_67_enex5;
  wire weight_write_data_data_and_68_enex5;
  wire weight_write_data_data_and_69_enex5;
  wire weight_write_data_data_and_70_enex5;
  wire weight_write_data_data_and_71_enex5;
  wire weight_write_data_data_and_72_enex5;
  wire weight_write_data_data_and_73_enex5;
  wire weight_write_data_data_and_74_enex5;
  wire weight_write_data_data_and_75_enex5;
  wire weight_write_data_data_and_76_enex5;
  wire weight_write_data_data_and_77_enex5;
  wire weight_write_data_data_and_78_enex5;
  wire weight_write_data_data_and_79_enex5;
  wire weight_write_addrs_and_2_enex5;
  wire weight_read_addrs_and_29_enex5;
  wire pe_config_UpdateManagerCounter_if_if_and_enex5;
  wire weight_port_read_out_data_and_244_enex5;
  wire weight_port_read_out_data_and_245_enex5;
  wire weight_port_read_out_data_and_246_enex5;
  wire PEManager_15U_PEManagerWrite_and_enex5;
  wire input_mem_banks_read_read_data_and_39_enex5;
  wire input_mem_banks_read_read_data_and_40_enex5;
  wire input_mem_banks_read_read_data_and_41_enex5;
  wire input_mem_banks_read_read_data_and_42_enex5;
  wire input_mem_banks_read_1_read_data_and_6_enex5;
  wire weight_read_addrs_and_30_enex5;
  wire rva_out_reg_data_and_143_enex5;
  wire rva_out_reg_data_and_144_enex5;
  wire rva_out_reg_data_and_145_enex5;
  wire weight_port_read_out_data_and_247_enex5;
  wire rva_out_reg_data_and_146_enex5;
  wire rva_out_reg_data_and_147_enex5;
  wire rva_out_reg_data_and_148_enex5;
  wire rva_out_reg_data_and_149_enex5;
  wire rva_out_reg_data_and_150_enex5;
  wire rva_out_reg_data_and_151_enex5;
  wire rva_out_reg_data_and_152_enex5;
  wire rva_out_reg_data_and_153_enex5;
  wire rva_out_reg_data_and_154_enex5;
  wire rva_out_reg_data_and_155_enex5;
  wire rva_out_reg_data_and_156_enex5;
  wire weight_mem_write_arbxbar_xbar_for_empty_and_enex5;
  wire input_mem_banks_read_read_data_and_43_enex5;
  wire input_mem_banks_read_read_data_and_44_enex5;
  wire input_mem_banks_read_read_data_and_45_enex5;
  wire input_mem_banks_read_read_data_and_46_enex5;
  wire input_mem_banks_read_1_read_data_and_7_enex5;
  wire rva_out_reg_data_and_157_enex5;
  wire rva_out_reg_data_and_158_enex5;
  wire rva_out_reg_data_and_159_enex5;
  wire rva_out_reg_data_and_160_enex5;
  wire rva_out_reg_data_and_161_enex5;
  wire rva_out_reg_data_and_162_enex5;
  wire rva_out_reg_data_and_163_enex5;
  wire rva_out_reg_data_and_164_enex5;
  wire rva_out_reg_data_and_165_enex5;
  wire rva_out_reg_data_and_166_enex5;
  wire rva_out_reg_data_and_167_enex5;
  wire input_mem_banks_read_read_data_and_33_enex5;
  wire rva_out_reg_data_and_168_enex5;
  wire rva_out_reg_data_and_169_enex5;
  wire rva_out_reg_data_and_170_enex5;
  wire rva_out_reg_data_and_171_enex5;
  wire rva_out_reg_data_and_172_enex5;
  wire rva_out_reg_data_and_173_enex5;
  wire rva_out_reg_data_and_174_enex5;
  wire rva_out_reg_data_and_175_enex5;
  wire input_mem_banks_read_read_data_and_34_enex5;
  wire rva_out_reg_data_and_176_enex5;
  wire rva_out_reg_data_and_177_enex5;
  wire rva_out_reg_data_and_178_enex5;
  wire rva_out_reg_data_and_179_enex5;
  wire rva_out_reg_data_and_180_enex5;
  wire rva_out_reg_data_and_181_enex5;
  wire rva_out_reg_data_and_117_enex5;
  wire rva_out_reg_data_and_182_enex5;
  wire rva_out_reg_data_and_183_enex5;
  wire rva_out_reg_data_and_184_enex5;
  wire rva_out_reg_data_and_185_enex5;
  wire rva_out_reg_data_and_186_enex5;
  wire weight_port_read_out_data_and_248_enex5;
  wire weight_port_read_out_data_and_249_enex5;
  wire weight_port_read_out_data_and_250_enex5;
  wire weight_port_read_out_data_and_251_enex5;
  wire weight_port_read_out_data_and_252_enex5;
  wire weight_port_read_out_data_and_253_enex5;
  wire weight_port_read_out_data_and_254_enex5;
  wire weight_port_read_out_data_and_255_enex5;
  wire weight_port_read_out_data_and_256_enex5;
  wire weight_port_read_out_data_and_257_enex5;
  wire weight_port_read_out_data_and_258_enex5;
  wire rva_out_reg_data_and_187_enex5;
  wire rva_out_reg_data_and_188_enex5;
  wire rva_out_reg_data_and_189_enex5;
  wire rva_out_reg_data_and_190_enex5;
  wire rva_out_reg_data_and_191_enex5;
  wire rva_out_reg_data_and_192_enex5;
  wire rva_out_reg_data_and_193_enex5;
  wire rva_out_reg_data_and_194_enex5;
  wire rva_out_reg_data_and_195_enex5;
  wire rva_out_reg_data_and_196_enex5;
  wire rva_out_reg_data_and_197_enex5;
  wire rva_out_reg_data_and_198_enex5;
  wire rva_out_reg_data_and_199_enex5;
  wire rva_out_reg_data_and_200_enex5;
  wire data_in_tmp_operator_2_for_and_15_tmp;
  wire data_in_tmp_operator_2_for_and_31_tmp;
  wire pe_manager_base_input_and_tmp;
  wire rva_in_reg_data_and_tmp;
  wire input_mem_banks_read_1_read_data_and_4_tmp;
  wire and_1434_tmp;
  wire and_1538_tmp;
  wire mux_433_itm;
  wire mux_47_itm;
  wire [30:0] accum_vector_data_acc_20_itm;
  wire [31:0] nl_accum_vector_data_acc_20_itm;
  wire [30:0] accum_vector_data_acc_14_itm;
  wire [31:0] nl_accum_vector_data_acc_14_itm;
  wire [30:0] accum_vector_data_acc_23_itm;
  wire [31:0] nl_accum_vector_data_acc_23_itm;
  wire [30:0] accum_vector_data_acc_11_itm;
  wire [31:0] nl_accum_vector_data_acc_11_itm;
  wire [30:0] accum_vector_data_acc_26_itm;
  wire [31:0] nl_accum_vector_data_acc_26_itm;
  wire [30:0] accum_vector_data_acc_8_itm;
  wire [31:0] nl_accum_vector_data_acc_8_itm;
  wire [30:0] accum_vector_data_acc_itm;
  wire [31:0] nl_accum_vector_data_acc_itm;
  wire [30:0] accum_vector_data_acc_17_itm;
  wire [31:0] nl_accum_vector_data_acc_17_itm;
  wire mux_260_itm;
  wire mux_258_itm;
  wire PECore_PushAxiRsp_if_else_mux_24_itm;
  wire PECore_PushAxiRsp_if_else_mux_25_itm;
  wire PECore_PushAxiRsp_if_else_mux_26_itm;
  wire mux_540_itm;
  wire accum_vector_data_and_55_cse;
  wire accum_vector_data_and_cse;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27;
  wire mux_101_nl;
  wire mux_100_nl;
  wire or_359_nl;
  wire or_358_nl;
  wire mux_104_nl;
  wire mux_103_nl;
  wire or_363_nl;
  wire or_362_nl;
  wire mux_107_nl;
  wire mux_106_nl;
  wire or_370_nl;
  wire or_369_nl;
  wire mux_110_nl;
  wire mux_109_nl;
  wire or_376_nl;
  wire or_836_nl;
  wire mux_114_nl;
  wire mux_113_nl;
  wire or_382_nl;
  wire or_837_nl;
  wire mux_117_nl;
  wire mux_116_nl;
  wire or_388_nl;
  wire or_838_nl;
  wire mux_120_nl;
  wire mux_119_nl;
  wire or_394_nl;
  wire or_839_nl;
  wire mux_124_nl;
  wire mux_123_nl;
  wire or_400_nl;
  wire or_399_nl;
  wire and_1075_nl;
  wire and_755_nl;
  wire mux_135_nl;
  wire mux_134_nl;
  wire mux_133_nl;
  wire and_759_nl;
  wire mux_129_nl;
  wire mux_132_nl;
  wire mux_131_nl;
  wire mux_130_nl;
  wire mux_428_nl;
  wire or_405_nl;
  wire or_404_nl;
  wire mux_138_nl;
  wire mux_137_nl;
  wire or_403_nl;
  wire or_402_nl;
  wire mux_437_nl;
  wire mux_436_nl;
  wire or_851_nl;
  wire mux_435_nl;
  wire nor_nl;
  wire PECore_UpdateFSM_switch_lp_not_23_nl;
  wire PECore_UpdateFSM_switch_lp_not_24_nl;
  wire PECore_UpdateFSM_switch_lp_not_25_nl;
  wire PECore_UpdateFSM_switch_lp_not_26_nl;
  wire PECore_UpdateFSM_switch_lp_not_27_nl;
  wire PECore_UpdateFSM_switch_lp_not_28_nl;
  wire PECore_UpdateFSM_switch_lp_not_29_nl;
  wire PECore_UpdateFSM_switch_lp_not_19_nl;
  wire accum_vector_operator_1_for_not_39_nl;
  wire accum_vector_operator_1_for_not_38_nl;
  wire accum_vector_operator_1_for_not_37_nl;
  wire accum_vector_operator_1_for_not_36_nl;
  wire accum_vector_operator_1_for_not_35_nl;
  wire accum_vector_operator_1_for_not_34_nl;
  wire[7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_1_nl;
  wire[7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl;
  wire weight_mem_run_3_for_5_and_177_nl;
  wire mux_460_nl;
  wire and_1270_nl;
  wire and_1269_nl;
  wire weight_mem_run_3_for_5_and_188_nl;
  wire weight_mem_run_3_for_5_and_191_nl;
  wire mux_462_nl;
  wire and_1275_nl;
  wire and_1274_nl;
  wire mux_18_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_136_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl;
  wire mux_21_nl;
  wire mux_20_nl;
  wire or_52_nl;
  wire mux_19_nl;
  wire or_50_nl;
  wire or_48_nl;
  wire mux_22_nl;
  wire nor_347_nl;
  wire mux_23_nl;
  wire mux_464_nl;
  wire mux_463_nl;
  wire nor_559_nl;
  wire nor_560_nl;
  wire[10:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl;
  wire[3:0] PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl;
  wire and_638_nl;
  wire[3:0] operator_4_false_acc_nl;
  wire[4:0] nl_operator_4_false_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_7_nl;
  wire mux_465_nl;
  wire mux_466_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_and_1_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_mux1h_18_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_nor_8_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_189_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_219_nl;
  wire mux_35_nl;
  wire mux_34_nl;
  wire or_196_nl;
  wire or_195_nl;
  wire or_194_nl;
  wire mux_467_nl;
  wire mux_486_nl;
  wire mux_485_nl;
  wire mux_36_nl;
  wire nor_350_nl;
  wire nand_39_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_134_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_151_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_28_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl;
  wire mux_490_nl;
  wire mux_489_nl;
  wire nor_584_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_48_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl;
  wire mux_37_nl;
  wire nor_355_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_80_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_138_nl;
  wire mux_38_nl;
  wire nor_356_nl;
  wire or_208_nl;
  wire mux_43_nl;
  wire mux_42_nl;
  wire nand_2_nl;
  wire mux_41_nl;
  wire nor_359_nl;
  wire mux_40_nl;
  wire or_225_nl;
  wire nor_360_nl;
  wire mux_39_nl;
  wire or_219_nl;
  wire or_217_nl;
  wire mux_592_nl;
  wire mux_60_nl;
  wire or_233_nl;
  wire mux_59_nl;
  wire mux_58_nl;
  wire mux_57_nl;
  wire mux_56_nl;
  wire mux_55_nl;
  wire mux_54_nl;
  wire mux_53_nl;
  wire mux_49_nl;
  wire mux_48_nl;
  wire mux_44_nl;
  wire or_228_nl;
  wire or_226_nl;
  wire mux_62_nl;
  wire mux_61_nl;
  wire nand_3_nl;
  wire or_236_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl;
  wire[7:0] PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_1_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_27_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_135_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_142_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_132_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_235_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_250_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_175_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_190_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_205_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_220_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_236_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_251_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_176_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_191_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_206_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_221_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_237_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_252_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_177_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_192_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_207_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_222_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_238_nl;
  wire mux_497_nl;
  wire mux_496_nl;
  wire nor_594_nl;
  wire mux_495_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_253_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_178_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_193_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_208_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_223_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_239_nl;
  wire mux_503_nl;
  wire mux_502_nl;
  wire nor_595_nl;
  wire mux_501_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_254_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_179_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_194_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_209_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_224_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_255_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_180_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_195_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_210_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_225_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_241_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_181_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_196_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_211_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_226_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_242_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_257_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_182_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_197_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_212_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_227_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_243_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_183_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_198_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_213_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_228_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_244_nl;
  wire mux_67_nl;
  wire mux_66_nl;
  wire nor_320_nl;
  wire[7:0] mux1h_6_nl;
  wire not_2283_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_199_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_229_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_245_nl;
  wire[7:0] mux1h_7_nl;
  wire not_2285_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_200_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_230_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_246_nl;
  wire[7:0] mux1h_8_nl;
  wire not_2287_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_201_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_231_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_247_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_202_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_232_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_248_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_203_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_233_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_140_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl;
  wire mux_73_nl;
  wire mux_74_nl;
  wire nor_371_nl;
  wire nor_16_nl;
  wire[7:0] input_mem_banks_read_1_for_mux_nl;
  wire and_1073_nl;
  wire mux_75_nl;
  wire or_829_nl;
  wire nor_373_nl;
  wire mux_81_nl;
  wire mux_80_nl;
  wire mux_79_nl;
  wire mux_78_nl;
  wire mux_77_nl;
  wire nor_379_nl;
  wire nor_380_nl;
  wire nor_381_nl;
  wire nor_382_nl;
  wire nor_383_nl;
  wire weight_port_read_out_data_mux_106_nl;
  wire and_667_nl;
  wire nor_499_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_234_nl;
  wire mux_82_nl;
  wire or_328_nl;
  wire or_327_nl;
  wire mux_90_nl;
  wire mux_89_nl;
  wire mux_88_nl;
  wire mux_86_nl;
  wire mux_85_nl;
  wire or_326_nl;
  wire mux_84_nl;
  wire mux_83_nl;
  wire mux_507_nl;
  wire mux_506_nl;
  wire mux_505_nl;
  wire or_1099_nl;
  wire mux_91_nl;
  wire mux_92_nl;
  wire[14:0] while_if_while_if_and_2_nl;
  wire mux_168_nl;
  wire or_511_nl;
  wire mux_167_nl;
  wire and_682_nl;
  wire or_512_nl;
  wire mux_94_nl;
  wire mux_93_nl;
  wire and_748_nl;
  wire or_334_nl;
  wire mux_95_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl;
  wire mux_96_nl;
  wire mux_97_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl;
  wire[30:0] accum_vector_data_acc_21_nl;
  wire[32:0] nl_accum_vector_data_acc_21_nl;
  wire[30:0] accum_vector_data_mux_57_nl;
  wire[30:0] accum_vector_data_mux_55_nl;
  wire[30:0] accum_vector_data_mux_53_nl;
  wire[30:0] accum_vector_data_acc_22_nl;
  wire[32:0] nl_accum_vector_data_acc_22_nl;
  wire[30:0] accum_vector_data_mux_51_nl;
  wire[30:0] accum_vector_data_mux_49_nl;
  wire[30:0] accum_vector_data_mux_47_nl;
  wire[30:0] accum_vector_data_acc_15_nl;
  wire[32:0] nl_accum_vector_data_acc_15_nl;
  wire[30:0] accum_vector_data_mux_79_nl;
  wire[30:0] accum_vector_data_mux_77_nl;
  wire[30:0] accum_vector_data_mux_75_nl;
  wire[30:0] accum_vector_data_acc_16_nl;
  wire[32:0] nl_accum_vector_data_acc_16_nl;
  wire[30:0] accum_vector_data_mux_73_nl;
  wire[30:0] accum_vector_data_mux_71_nl;
  wire[30:0] accum_vector_data_mux_69_nl;
  wire[30:0] accum_vector_data_acc_24_nl;
  wire[32:0] nl_accum_vector_data_acc_24_nl;
  wire[30:0] accum_vector_data_mux_45_nl;
  wire[30:0] accum_vector_data_mux_43_nl;
  wire[30:0] accum_vector_data_mux_41_nl;
  wire[30:0] accum_vector_data_acc_25_nl;
  wire[32:0] nl_accum_vector_data_acc_25_nl;
  wire[30:0] accum_vector_data_mux_39_nl;
  wire[30:0] accum_vector_data_mux_37_nl;
  wire[30:0] accum_vector_data_acc_12_nl;
  wire[32:0] nl_accum_vector_data_acc_12_nl;
  wire[30:0] accum_vector_data_mux_89_nl;
  wire[30:0] accum_vector_data_mux_87_nl;
  wire[30:0] accum_vector_data_mux_85_nl;
  wire[30:0] accum_vector_data_acc_13_nl;
  wire[32:0] nl_accum_vector_data_acc_13_nl;
  wire[30:0] accum_vector_data_mux_83_nl;
  wire[30:0] accum_vector_data_mux_81_nl;
  wire[30:0] accum_vector_data_acc_27_nl;
  wire[32:0] nl_accum_vector_data_acc_27_nl;
  wire[30:0] accum_vector_data_mux_35_nl;
  wire[30:0] accum_vector_data_mux_33_nl;
  wire[30:0] accum_vector_data_mux_31_nl;
  wire[30:0] accum_vector_data_acc_28_nl;
  wire[32:0] nl_accum_vector_data_acc_28_nl;
  wire[30:0] accum_vector_data_mux_29_nl;
  wire[30:0] accum_vector_data_mux_27_nl;
  wire[30:0] accum_vector_data_acc_9_nl;
  wire[32:0] nl_accum_vector_data_acc_9_nl;
  wire[30:0] accum_vector_data_mux_99_nl;
  wire[30:0] accum_vector_data_mux_97_nl;
  wire[30:0] accum_vector_data_mux_95_nl;
  wire[30:0] accum_vector_data_acc_10_nl;
  wire[32:0] nl_accum_vector_data_acc_10_nl;
  wire[30:0] accum_vector_data_mux_93_nl;
  wire[30:0] accum_vector_data_mux_91_nl;
  wire[30:0] accum_vector_data_acc_29_nl;
  wire[32:0] nl_accum_vector_data_acc_29_nl;
  wire[30:0] accum_vector_data_mux_25_nl;
  wire[30:0] accum_vector_data_mux_23_nl;
  wire[30:0] accum_vector_data_mux_21_nl;
  wire[30:0] accum_vector_data_acc_30_nl;
  wire[32:0] nl_accum_vector_data_acc_30_nl;
  wire[30:0] accum_vector_data_mux_19_nl;
  wire[30:0] accum_vector_data_mux_17_nl;
  wire[30:0] accum_vector_data_acc_18_nl;
  wire[32:0] nl_accum_vector_data_acc_18_nl;
  wire[30:0] accum_vector_data_mux_67_nl;
  wire[30:0] accum_vector_data_mux_65_nl;
  wire[30:0] accum_vector_data_mux_63_nl;
  wire[30:0] accum_vector_data_acc_19_nl;
  wire[32:0] nl_accum_vector_data_acc_19_nl;
  wire[30:0] accum_vector_data_mux_61_nl;
  wire[30:0] accum_vector_data_mux_59_nl;
  wire[30:0] ProductSum_for_mux_nl;
  wire accum_vector_operator_1_for_not_56_nl;
  wire[30:0] ProductSum_for_mux_1_nl;
  wire accum_vector_operator_1_for_not_57_nl;
  wire[30:0] ProductSum_for_mux_2_nl;
  wire accum_vector_operator_1_for_not_58_nl;
  wire[30:0] ProductSum_for_mux_3_nl;
  wire accum_vector_operator_1_for_not_59_nl;
  wire[30:0] ProductSum_for_mux_4_nl;
  wire accum_vector_operator_1_for_not_40_nl;
  wire[30:0] ProductSum_for_mux_5_nl;
  wire accum_vector_operator_1_for_not_60_nl;
  wire[30:0] ProductSum_for_mux_6_nl;
  wire accum_vector_operator_1_for_not_61_nl;
  wire[30:0] ProductSum_for_mux_7_nl;
  wire accum_vector_operator_1_for_not_62_nl;
  wire[30:0] ProductSum_for_mux_8_nl;
  wire accum_vector_operator_1_for_not_63_nl;
  wire[30:0] ProductSum_for_mux_9_nl;
  wire accum_vector_operator_1_for_not_42_nl;
  wire[30:0] ProductSum_for_mux_10_nl;
  wire accum_vector_operator_1_for_not_64_nl;
  wire[30:0] ProductSum_for_mux_11_nl;
  wire accum_vector_operator_1_for_not_65_nl;
  wire[30:0] ProductSum_for_mux_12_nl;
  wire accum_vector_operator_1_for_not_66_nl;
  wire[30:0] ProductSum_for_mux_13_nl;
  wire accum_vector_operator_1_for_not_67_nl;
  wire[30:0] ProductSum_for_mux_14_nl;
  wire accum_vector_operator_1_for_not_44_nl;
  wire[30:0] ProductSum_for_mux_15_nl;
  wire accum_vector_operator_1_for_not_68_nl;
  wire[30:0] ProductSum_for_mux_16_nl;
  wire accum_vector_operator_1_for_not_69_nl;
  wire[30:0] ProductSum_for_mux_17_nl;
  wire accum_vector_operator_1_for_not_70_nl;
  wire[30:0] ProductSum_for_mux_18_nl;
  wire accum_vector_operator_1_for_not_71_nl;
  wire[30:0] ProductSum_for_mux_19_nl;
  wire accum_vector_operator_1_for_not_72_nl;
  wire[30:0] ProductSum_for_mux_20_nl;
  wire accum_vector_operator_1_for_not_46_nl;
  wire[30:0] ProductSum_for_mux_21_nl;
  wire accum_vector_operator_1_for_not_73_nl;
  wire[30:0] ProductSum_for_mux_22_nl;
  wire accum_vector_operator_1_for_not_74_nl;
  wire[30:0] ProductSum_for_mux_23_nl;
  wire accum_vector_operator_1_for_not_75_nl;
  wire[30:0] ProductSum_for_mux_24_nl;
  wire accum_vector_operator_1_for_not_76_nl;
  wire[30:0] ProductSum_for_mux_25_nl;
  wire accum_vector_operator_1_for_not_48_nl;
  wire[30:0] ProductSum_for_mux_26_nl;
  wire accum_vector_operator_1_for_not_77_nl;
  wire[30:0] ProductSum_for_mux_27_nl;
  wire accum_vector_operator_1_for_not_78_nl;
  wire[30:0] ProductSum_for_mux_28_nl;
  wire accum_vector_operator_1_for_not_79_nl;
  wire[30:0] ProductSum_for_mux_29_nl;
  wire accum_vector_operator_1_for_not_80_nl;
  wire[30:0] ProductSum_for_mux_30_nl;
  wire accum_vector_operator_1_for_not_81_nl;
  wire[30:0] ProductSum_for_mux_31_nl;
  wire accum_vector_operator_1_for_not_50_nl;
  wire[30:0] ProductSum_for_mux_32_nl;
  wire accum_vector_operator_1_for_not_82_nl;
  wire[30:0] ProductSum_for_mux_33_nl;
  wire accum_vector_operator_1_for_not_83_nl;
  wire[30:0] ProductSum_for_mux_34_nl;
  wire accum_vector_operator_1_for_not_84_nl;
  wire[30:0] ProductSum_for_mux_35_nl;
  wire accum_vector_operator_1_for_not_85_nl;
  wire[30:0] ProductSum_for_mux_36_nl;
  wire accum_vector_operator_1_for_not_52_nl;
  wire[30:0] ProductSum_for_mux_37_nl;
  wire accum_vector_operator_1_for_not_86_nl;
  wire[30:0] ProductSum_for_mux_38_nl;
  wire accum_vector_operator_1_for_not_87_nl;
  wire[30:0] ProductSum_for_mux_39_nl;
  wire accum_vector_operator_1_for_not_88_nl;
  wire[30:0] ProductSum_for_mux_40_nl;
  wire accum_vector_operator_1_for_not_89_nl;
  wire[30:0] ProductSum_for_mux_41_nl;
  wire accum_vector_operator_1_for_not_54_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_56_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_57_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_58_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_59_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_60_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_61_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_74_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_84_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_85_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl;
  wire[14:0] PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_nl;
  wire[14:0] nl_operator_15_false_acc_nl;
  wire[14:0] PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[12:0] operator_15_false_acc_1_nl;
  wire[13:0] nl_operator_15_false_acc_1_nl;
  wire[14:0] PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_2_nl;
  wire[14:0] nl_operator_15_false_acc_2_nl;
  wire[14:0] PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl;
  wire[7:0] pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl;
  wire[7:0] operator_8_false_acc_nl;
  wire[8:0] nl_operator_8_false_acc_nl;
  wire pe_config_UpdateInputCounter_not_nl;
  wire pe_config_input_counter_nand_nl;
  wire[7:0] pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl;
  wire[7:0] operator_8_false_1_acc_nl;
  wire[8:0] nl_operator_8_false_1_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_9_nl;
  wire pe_config_output_counter_nand_nl;
  wire while_and_152_nl;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl;
  wire while_if_or_nl;
  wire while_if_and_4_nl;
  wire[7:0] mux1h_11_nl;
  wire not_2293_nl;
  wire[7:0] mux1h_12_nl;
  wire and_1066_nl;
  wire and_1067_nl;
  wire and_1068_nl;
  wire and_1069_nl;
  wire and_1070_nl;
  wire and_1071_nl;
  wire nor_512_nl;
  wire not_2295_nl;
  wire PECore_PushAxiRsp_mux_25_nl;
  wire[7:0] while_if_while_if_and_27_nl;
  wire[7:0] while_if_while_if_and_28_nl;
  wire[7:0] while_if_while_if_and_30_nl;
  wire[7:0] while_if_while_if_and_31_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_220_nl;
  wire or_565_nl;
  wire mux_219_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_256_nl;
  wire mux_255_nl;
  wire mux_254_nl;
  wire or_612_nl;
  wire or_607_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl;
  wire mux_287_nl;
  wire nor_500_nl;
  wire nor_501_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl;
  wire nor_502_nl;
  wire mux_323_nl;
  wire mux_322_nl;
  wire mux_321_nl;
  wire or_708_nl;
  wire or_706_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_24_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl;
  wire and_709_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_360_nl;
  wire mux_359_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl;
  wire mux_398_nl;
  wire nor_503_nl;
  wire nor_504_nl;
  wire mux_397_nl;
  wire mux_396_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_44_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_46_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_47_nl;
  wire PECore_UpdateFSM_switch_lp_mux1h_14_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl;
  wire PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl;
  wire PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_nl;
  wire weight_mem_banks_load_store_1_for_else_else_or_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_4_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_6_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_8_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_265_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_21_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_108_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_148_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_124_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_163_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_107_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_149_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_123_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_164_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_102_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_151_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_118_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_166_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_105_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_152_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_121_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_167_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_104_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_153_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_120_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_168_nl;
  wire[7:0] PEManager_15U_GetInputAddr_acc_nl;
  wire[8:0] nl_PEManager_15U_GetInputAddr_acc_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_589_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_590_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_591_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_592_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_593_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_594_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_595_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_596_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_597_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_598_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_599_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_600_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_603_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_604_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_605_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_606_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_607_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_608_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_609_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_619_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_620_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_621_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_622_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_624_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_627_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_628_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_630_nl;
  wire or_36_nl;
  wire mux_28_nl;
  wire mux_27_nl;
  wire mux_26_nl;
  wire and_735_nl;
  wire or_230_nl;
  wire or_232_nl;
  wire mux_51_nl;
  wire mux_99_nl;
  wire or_357_nl;
  wire mux_102_nl;
  wire or_361_nl;
  wire mux_105_nl;
  wire or_365_nl;
  wire mux_108_nl;
  wire or_373_nl;
  wire or_381_nl;
  wire or_380_nl;
  wire mux_112_nl;
  wire or_379_nl;
  wire mux_115_nl;
  wire or_385_nl;
  wire mux_118_nl;
  wire or_391_nl;
  wire or_398_nl;
  wire or_397_nl;
  wire mux_122_nl;
  wire or_396_nl;
  wire mux_160_nl;
  wire or_494_nl;
  wire mux_159_nl;
  wire or_493_nl;
  wire nor_35_nl;
  wire or_513_nl;
  wire or_518_nl;
  wire mux_173_nl;
  wire mux_172_nl;
  wire mux_171_nl;
  wire or_517_nl;
  wire or_515_nl;
  wire mux_179_nl;
  wire mux_178_nl;
  wire mux_177_nl;
  wire mux_176_nl;
  wire mux_175_nl;
  wire or_522_nl;
  wire or_520_nl;
  wire mux_184_nl;
  wire mux_183_nl;
  wire mux_182_nl;
  wire nand_9_nl;
  wire mux_189_nl;
  wire mux_188_nl;
  wire mux_187_nl;
  wire or_526_nl;
  wire mux_186_nl;
  wire or_525_nl;
  wire or_523_nl;
  wire mux_191_nl;
  wire or_527_nl;
  wire mux_194_nl;
  wire or_537_nl;
  wire or_538_nl;
  wire or_533_nl;
  wire mux_200_nl;
  wire or_541_nl;
  wire mux_199_nl;
  wire or_539_nl;
  wire mux_208_nl;
  wire mux_207_nl;
  wire or_551_nl;
  wire mux_206_nl;
  wire mux_205_nl;
  wire mux_204_nl;
  wire mux_203_nl;
  wire or_550_nl;
  wire mux_202_nl;
  wire or_547_nl;
  wire mux_201_nl;
  wire or_546_nl;
  wire or_545_nl;
  wire mux_211_nl;
  wire mux_210_nl;
  wire or_557_nl;
  wire or_556_nl;
  wire or_555_nl;
  wire or_554_nl;
  wire mux_218_nl;
  wire mux_217_nl;
  wire mux_216_nl;
  wire mux_215_nl;
  wire mux_214_nl;
  wire mux_213_nl;
  wire or_564_nl;
  wire or_563_nl;
  wire or_562_nl;
  wire or_561_nl;
  wire or_558_nl;
  wire mux_222_nl;
  wire mux_221_nl;
  wire or_569_nl;
  wire or_567_nl;
  wire mux_225_nl;
  wire mux_224_nl;
  wire nand_10_nl;
  wire mux_228_nl;
  wire mux_227_nl;
  wire nand_11_nl;
  wire mux_231_nl;
  wire mux_230_nl;
  wire or_571_nl;
  wire or_570_nl;
  wire mux_235_nl;
  wire mux_234_nl;
  wire mux_233_nl;
  wire or_576_nl;
  wire or_575_nl;
  wire or_574_nl;
  wire mux_239_nl;
  wire mux_238_nl;
  wire mux_237_nl;
  wire or_583_nl;
  wire or_582_nl;
  wire mux_245_nl;
  wire mux_244_nl;
  wire mux_243_nl;
  wire or_590_nl;
  wire or_589_nl;
  wire mux_242_nl;
  wire mux_241_nl;
  wire or_588_nl;
  wire or_587_nl;
  wire mux_240_nl;
  wire or_586_nl;
  wire or_579_nl;
  wire mux_253_nl;
  wire mux_252_nl;
  wire mux_251_nl;
  wire mux_250_nl;
  wire nor_432_nl;
  wire nor_433_nl;
  wire nor_434_nl;
  wire nor_435_nl;
  wire mux_249_nl;
  wire mux_248_nl;
  wire mux_247_nl;
  wire nor_436_nl;
  wire nor_437_nl;
  wire nor_438_nl;
  wire nor_439_nl;
  wire nand_13_nl;
  wire nand_12_nl;
  wire mux_271_nl;
  wire mux_270_nl;
  wire mux_269_nl;
  wire mux_268_nl;
  wire mux_267_nl;
  wire mux_266_nl;
  wire mux_265_nl;
  wire mux_264_nl;
  wire mux_263_nl;
  wire mux_262_nl;
  wire mux_261_nl;
  wire or_620_nl;
  wire mux_259_nl;
  wire or_617_nl;
  wire nor_441_nl;
  wire mux_278_nl;
  wire mux_277_nl;
  wire or_635_nl;
  wire mux_276_nl;
  wire or_634_nl;
  wire or_633_nl;
  wire nor_442_nl;
  wire mux_275_nl;
  wire mux_274_nl;
  wire or_627_nl;
  wire mux_273_nl;
  wire or_626_nl;
  wire or_625_nl;
  wire mux_286_nl;
  wire mux_285_nl;
  wire mux_284_nl;
  wire mux_283_nl;
  wire nor_443_nl;
  wire nor_444_nl;
  wire nor_445_nl;
  wire nor_446_nl;
  wire mux_282_nl;
  wire mux_281_nl;
  wire mux_280_nl;
  wire nor_447_nl;
  wire nor_448_nl;
  wire nor_449_nl;
  wire nor_450_nl;
  wire mux_290_nl;
  wire mux_289_nl;
  wire mux_288_nl;
  wire mux_292_nl;
  wire or_668_nl;
  wire mux_291_nl;
  wire or_664_nl;
  wire mux_296_nl;
  wire mux_295_nl;
  wire mux_294_nl;
  wire or_675_nl;
  wire or_670_nl;
  wire mux_298_nl;
  wire mux_297_nl;
  wire mux_302_nl;
  wire mux_301_nl;
  wire mux_307_nl;
  wire mux_306_nl;
  wire mux_305_nl;
  wire mux_304_nl;
  wire or_692_nl;
  wire mux_303_nl;
  wire or_690_nl;
  wire mux_300_nl;
  wire mux_299_nl;
  wire or_685_nl;
  wire or_684_nl;
  wire or_682_nl;
  wire mux_308_nl;
  wire or_696_nl;
  wire or_695_nl;
  wire or_700_nl;
  wire mux_311_nl;
  wire or_833_nl;
  wire or_699_nl;
  wire mux_320_nl;
  wire mux_319_nl;
  wire mux_318_nl;
  wire mux_317_nl;
  wire or_704_nl;
  wire or_703_nl;
  wire mux_316_nl;
  wire or_702_nl;
  wire or_701_nl;
  wire mux_315_nl;
  wire mux_314_nl;
  wire mux_313_nl;
  wire or_698_nl;
  wire or_694_nl;
  wire or_716_nl;
  wire or_713_nl;
  wire while_mux_1419_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_610_nl;
  wire mux_325_nl;
  wire mux_332_nl;
  wire mux_331_nl;
  wire mux_330_nl;
  wire mux_329_nl;
  wire or_723_nl;
  wire or_722_nl;
  wire or_721_nl;
  wire mux_328_nl;
  wire mux_327_nl;
  wire or_720_nl;
  wire or_719_nl;
  wire or_718_nl;
  wire or_725_nl;
  wire or_724_nl;
  wire mux_335_nl;
  wire mux_334_nl;
  wire or_728_nl;
  wire or_726_nl;
  wire or_735_nl;
  wire or_733_nl;
  wire mux_339_nl;
  wire mux_338_nl;
  wire or_742_nl;
  wire or_736_nl;
  wire or_746_nl;
  wire or_744_nl;
  wire or_750_nl;
  wire or_747_nl;
  wire mux_350_nl;
  wire mux_349_nl;
  wire mux_348_nl;
  wire nand_18_nl;
  wire or_756_nl;
  wire or_755_nl;
  wire mux_347_nl;
  wire mux_346_nl;
  wire mux_345_nl;
  wire or_754_nl;
  wire or_753_nl;
  wire mux_344_nl;
  wire mux_343_nl;
  wire or_752_nl;
  wire or_751_nl;
  wire mux_358_nl;
  wire mux_357_nl;
  wire mux_356_nl;
  wire mux_355_nl;
  wire nor_463_nl;
  wire nor_464_nl;
  wire nor_465_nl;
  wire nor_466_nl;
  wire mux_354_nl;
  wire mux_353_nl;
  wire mux_352_nl;
  wire nor_467_nl;
  wire nor_468_nl;
  wire nor_469_nl;
  wire nor_470_nl;
  wire or_769_nl;
  wire or_768_nl;
  wire mux_365_nl;
  wire mux_364_nl;
  wire or_770_nl;
  wire or_767_nl;
  wire nand_19_nl;
  wire nand_20_nl;
  wire mux_377_nl;
  wire mux_376_nl;
  wire or_775_nl;
  wire mux_375_nl;
  wire nand_21_nl;
  wire mux_374_nl;
  wire mux_373_nl;
  wire mux_372_nl;
  wire mux_371_nl;
  wire mux_370_nl;
  wire or_774_nl;
  wire or_773_nl;
  wire or_781_nl;
  wire or_778_nl;
  wire nor_471_nl;
  wire mux_387_nl;
  wire or_794_nl;
  wire mux_386_nl;
  wire mux_385_nl;
  wire or_792_nl;
  wire or_791_nl;
  wire nor_472_nl;
  wire mux_384_nl;
  wire mux_383_nl;
  wire or_786_nl;
  wire mux_382_nl;
  wire or_784_nl;
  wire mux_381_nl;
  wire mux_395_nl;
  wire mux_394_nl;
  wire mux_393_nl;
  wire mux_392_nl;
  wire nor_473_nl;
  wire nor_474_nl;
  wire nor_475_nl;
  wire nor_476_nl;
  wire mux_391_nl;
  wire mux_390_nl;
  wire mux_389_nl;
  wire nor_477_nl;
  wire nor_478_nl;
  wire nor_479_nl;
  wire nor_480_nl;
  wire and_552_nl;
  wire and_550_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl;
  wire weight_mem_banks_write_if_for_if_and_35_nl;
  wire weight_mem_banks_write_if_for_if_and_36_nl;
  wire weight_mem_banks_write_if_for_if_and_37_nl;
  wire weight_mem_banks_write_if_for_if_and_38_nl;
  wire weight_mem_banks_write_if_for_if_and_39_nl;
  wire weight_mem_banks_write_if_for_if_and_40_nl;
  wire weight_mem_banks_write_if_for_if_and_41_nl;
  wire weight_mem_banks_write_if_for_if_mux_7_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl;
  wire mux_146_nl;
  wire nor_497_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl;
  wire weight_mem_banks_write_if_for_if_and_28_nl;
  wire weight_mem_banks_write_if_for_if_and_29_nl;
  wire weight_mem_banks_write_if_for_if_and_30_nl;
  wire weight_mem_banks_write_if_for_if_and_31_nl;
  wire weight_mem_banks_write_if_for_if_and_32_nl;
  wire weight_mem_banks_write_if_for_if_and_33_nl;
  wire weight_mem_banks_write_if_for_if_and_34_nl;
  wire weight_mem_banks_write_if_for_if_mux_6_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl;
  wire mux_145_nl;
  wire nor_496_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl;
  wire weight_mem_banks_write_if_for_if_and_21_nl;
  wire weight_mem_banks_write_if_for_if_and_22_nl;
  wire weight_mem_banks_write_if_for_if_and_23_nl;
  wire weight_mem_banks_write_if_for_if_and_24_nl;
  wire weight_mem_banks_write_if_for_if_and_25_nl;
  wire weight_mem_banks_write_if_for_if_and_26_nl;
  wire weight_mem_banks_write_if_for_if_and_27_nl;
  wire weight_mem_banks_write_if_for_if_mux_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl;
  wire mux_144_nl;
  wire nor_495_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl;
  wire weight_mem_banks_write_if_for_if_and_14_nl;
  wire weight_mem_banks_write_if_for_if_and_15_nl;
  wire weight_mem_banks_write_if_for_if_and_16_nl;
  wire weight_mem_banks_write_if_for_if_and_17_nl;
  wire weight_mem_banks_write_if_for_if_and_18_nl;
  wire weight_mem_banks_write_if_for_if_and_19_nl;
  wire weight_mem_banks_write_if_for_if_and_20_nl;
  wire weight_mem_banks_write_if_for_if_mux_4_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl;
  wire mux_143_nl;
  wire nor_494_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl;
  wire weight_mem_banks_write_if_for_if_and_7_nl;
  wire weight_mem_banks_write_if_for_if_and_8_nl;
  wire weight_mem_banks_write_if_for_if_and_9_nl;
  wire weight_mem_banks_write_if_for_if_and_10_nl;
  wire weight_mem_banks_write_if_for_if_and_11_nl;
  wire weight_mem_banks_write_if_for_if_and_12_nl;
  wire weight_mem_banks_write_if_for_if_and_13_nl;
  wire weight_mem_banks_write_if_for_if_mux_3_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl;
  wire mux_142_nl;
  wire nor_493_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl;
  wire weight_mem_banks_write_if_for_if_and_nl;
  wire weight_mem_banks_write_if_for_if_and_1_nl;
  wire weight_mem_banks_write_if_for_if_and_2_nl;
  wire weight_mem_banks_write_if_for_if_and_3_nl;
  wire weight_mem_banks_write_if_for_if_and_4_nl;
  wire weight_mem_banks_write_if_for_if_and_5_nl;
  wire weight_mem_banks_write_if_for_if_and_6_nl;
  wire weight_mem_banks_write_if_for_if_mux_2_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl;
  wire mux_141_nl;
  wire nor_492_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_1_nl;
  wire weight_mem_banks_write_if_for_if_mux_54_nl;
  wire mux_140_nl;
  wire nor_491_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_nl;
  wire weight_mem_banks_write_if_for_if_mux_53_nl;
  wire mux_139_nl;
  wire nor_490_nl;
  wire rva_out_reg_data_mux_37_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_23_nl;
  wire rva_out_reg_data_mux_38_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_24_nl;
  wire rva_out_reg_data_mux_39_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_25_nl;
  wire PECore_PushAxiRsp_if_else_mux_27_nl;
  wire rva_out_reg_data_mux_41_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_26_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_mux_22_nl;
  wire PECore_PushAxiRsp_if_else_mux_28_nl;
  wire rva_out_reg_data_mux_40_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl;
  wire mux_11_nl;
  wire mux_10_nl;
  wire mux_13_nl;
  wire mux_12_nl;
  wire nor_279_nl;
  wire mux_525_nl;
  wire mux_524_nl;
  wire mux_523_nl;
  wire[3:0] mux1h_3_nl;
  wire not_2368_nl;
  wire[3:0] mux1h_15_nl;
  wire not_2277_nl;
  wire mux1h_4_nl;
  wire[6:0] mux1h_13_nl;
  wire not_2366_nl;
  wire mux1h_5_nl;
  wire[6:0] mux1h_14_nl;
  wire not_2367_nl;
  wire mux_33_nl;
  wire mux_32_nl;
  wire mux_31_nl;
  wire mux_30_nl;
  wire mux_29_nl;
  wire or_191_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_3_nl;
  wire not_2269_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_87_nl;
  wire not_2270_nl;
  wire mux_64_nl;
  wire nor_319_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_76_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_88_nl;
  wire not_2272_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_81_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_89_nl;
  wire not_2274_nl;
  wire mux_72_nl;
  wire or_271_nl;
  wire mux_71_nl;
  wire nor_368_nl;
  wire nor_369_nl;
  wire mux_70_nl;
  wire mux_69_nl;
  wire mux_68_nl;
  wire or_263_nl;
  wire[3:0] mux_415_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_or_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_86_nl;
  wire not_2275_nl;
  wire[3:0] mux_416_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_or_1_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_90_nl;
  wire and_662_nl;
  wire not_2276_nl;
  wire[3:0] mux1h_9_nl;
  wire not_2369_nl;
  wire[3:0] mux1h_16_nl;
  wire not_2289_nl;
  wire[1:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_111_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_264_nl;
  wire[1:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_127_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_265_nl;
  wire[5:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_128_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_145_nl;
  wire[5:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_129_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_160_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_110_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_126_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_130_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_131_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_267_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_109_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_125_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_132_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_133_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_269_nl;
  wire mux_14_nl;
  wire or_33_nl;
  wire mux_545_nl;
  wire and_1544_nl;
  wire and_1543_nl;
  wire mux_547_nl;
  wire and_1549_nl;
  wire and_1548_nl;
  wire mux_554_nl;
  wire mux_553_nl;
  wire nor_616_nl;
  wire mux_552_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_134_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_240_nl;
  wire mux_564_nl;
  wire or_1179_nl;
  wire or_1177_nl;
  wire mux_563_nl;
  wire mux_562_nl;
  wire or_1176_nl;
  wire or_1175_nl;
  wire or_1174_nl;
  wire mux_76_nl;
  wire[5:0] while_if_while_if_and_35_nl;
  wire[6:0] while_if_while_if_and_34_nl;
  wire[6:0] while_if_while_if_and_33_nl;
  wire mux_581_nl;
  wire and_1579_nl;
  wire and_1578_nl;
  wire[3:0] mux1h_10_nl;
  wire not_2374_nl;
  wire[3:0] mux1h_17_nl;
  wire not_2291_nl;
  wire[3:0] while_if_while_if_and_29_nl;
  wire[3:0] while_if_while_if_and_36_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_106_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_271_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_122_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_272_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_135_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_150_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_136_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_165_nl;
  wire[3:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl;
  wire[3:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl;
  wire[3:0] PECore_DecodeAxiRead_switch_lp_mux_20_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_27_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_21_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_mux_28_nl;
  wire or_929_nl;
  wire or_933_nl;
  wire or_1054_nl;
  wire mux_493_nl;
  wire mux_492_nl;
  wire mux_521_nl;
  wire mux_520_nl;
  wire or_1122_nl;
  wire or_1121_nl;
  wire or_1120_nl;
  wire or_1125_nl;
  wire mux_539_nl;
  wire mux_538_nl;
  wire or_1146_nl;
  wire or_1145_nl;
  wire or_1144_nl;
  wire or_1149_nl;
  wire or_1151_nl;
  wire or_1155_nl;
  wire and_1626_nl;
  wire mux_550_nl;
  wire and_1627_nl;
  wire mux_549_nl;
  wire mux_548_nl;
  wire and_1628_nl;
  wire and_1629_nl;
  wire and_1630_nl;
  wire or_1204_nl;
  wire mux_491_nl;
  wire or_1051_nl;
  wire mux_543_nl;
  wire mux_542_nl;
  wire mux_541_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [30:0] nl_PECore_RunScale_if_for_4_mul_1_cmp_b;
  assign nl_PECore_RunScale_if_for_4_mul_1_cmp_b = MUX_v_31_2_2(accum_vector_data_3_sva,
      accum_vector_data_acc_17_itm, accum_vector_data_and_55_cse);
  wire [30:0] nl_PECore_RunScale_if_for_4_mul_1_cmp_1_b;
  assign nl_PECore_RunScale_if_for_4_mul_1_cmp_1_b = MUX_v_31_2_2(accum_vector_data_7_sva,
      accum_vector_data_acc_itm, accum_vector_data_and_55_cse);
  wire [30:0] nl_PECore_RunScale_if_for_4_mul_1_cmp_2_b;
  assign nl_PECore_RunScale_if_for_4_mul_1_cmp_2_b = MUX_v_31_2_2(accum_vector_data_0_sva,
      accum_vector_data_acc_8_itm, accum_vector_data_and_55_cse);
  wire [30:0] nl_PECore_RunScale_if_for_4_mul_1_cmp_3_b;
  assign nl_PECore_RunScale_if_for_4_mul_1_cmp_3_b = MUX_v_31_2_2(accum_vector_data_6_sva,
      accum_vector_data_acc_26_itm, accum_vector_data_and_55_cse);
  wire [30:0] nl_PECore_RunScale_if_for_4_mul_1_cmp_4_b;
  assign nl_PECore_RunScale_if_for_4_mul_1_cmp_4_b = MUX_v_31_2_2(accum_vector_data_1_sva,
      accum_vector_data_acc_11_itm, accum_vector_data_and_55_cse);
  wire [30:0] nl_PECore_RunScale_if_for_4_mul_1_cmp_5_b;
  assign nl_PECore_RunScale_if_for_4_mul_1_cmp_5_b = MUX_v_31_2_2(accum_vector_data_5_sva,
      accum_vector_data_acc_23_itm, accum_vector_data_and_55_cse);
  wire [30:0] nl_PECore_RunScale_if_for_4_mul_1_cmp_6_b;
  assign nl_PECore_RunScale_if_for_4_mul_1_cmp_6_b = MUX_v_31_2_2(accum_vector_data_2_sva,
      accum_vector_data_acc_14_itm, accum_vector_data_and_55_cse);
  wire [30:0] nl_PECore_RunScale_if_for_4_mul_1_cmp_7_b;
  assign nl_PECore_RunScale_if_for_4_mul_1_cmp_7_b = MUX_v_31_2_2(accum_vector_data_4_sva,
      accum_vector_data_acc_20_itm, accum_vector_data_and_55_cse);
  wire  nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (~ reg_rva_in_reg_rw_sva_2_cse);
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0];
  wire  nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a = PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2
      & reg_rva_in_reg_rw_sva_2_cse;
  wire [2:0] nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s = weight_write_addrs_lpi_1_dfm_1_2[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s = {(weight_read_addrs_6_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_4[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s = weight_read_addrs_7_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s = {(weight_read_addrs_2_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s = {(weight_read_addrs_4_14_2_lpi_1_dfm_1_1[0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[1:0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s = weight_read_addrs_3_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s = weight_read_addrs_5_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s = weight_read_addrs_1_lpi_1_dfm_1_1[2:0];
  wire[27:0] act_port_reg_data_mux_7_nl;
  wire[27:0] act_port_reg_data_mux_6_nl;
  wire[27:0] act_port_reg_data_mux_5_nl;
  wire[27:0] act_port_reg_data_mux_4_nl;
  wire[27:0] act_port_reg_data_mux_3_nl;
  wire[27:0] act_port_reg_data_mux_2_nl;
  wire[27:0] act_port_reg_data_mux_1_nl;
  wire[27:0] act_port_reg_data_mux_nl;
  wire [255:0] nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign act_port_reg_data_mux_7_nl = MUX_v_28_2_2(act_port_reg_data_251_224_sva,
      (PECore_RunScale_if_for_4_mul_1_cmp_1_z[38:11]), act_port_reg_data_and_16_cse);
  assign act_port_reg_data_mux_6_nl = MUX_v_28_2_2(act_port_reg_data_219_192_sva,
      (PECore_RunScale_if_for_4_mul_1_cmp_3_z[38:11]), act_port_reg_data_and_16_cse);
  assign act_port_reg_data_mux_5_nl = MUX_v_28_2_2(act_port_reg_data_187_160_sva,
      (PECore_RunScale_if_for_4_mul_1_cmp_5_z[38:11]), act_port_reg_data_and_16_cse);
  assign act_port_reg_data_mux_4_nl = MUX_v_28_2_2(act_port_reg_data_155_128_sva,
      (PECore_RunScale_if_for_4_mul_1_cmp_7_z[38:11]), act_port_reg_data_and_16_cse);
  assign act_port_reg_data_mux_3_nl = MUX_v_28_2_2(act_port_reg_data_123_96_sva,
      (PECore_RunScale_if_for_4_mul_1_cmp_z[38:11]), act_port_reg_data_and_16_cse);
  assign act_port_reg_data_mux_2_nl = MUX_v_28_2_2(act_port_reg_data_91_64_sva, (PECore_RunScale_if_for_4_mul_1_cmp_6_z[38:11]),
      act_port_reg_data_and_16_cse);
  assign act_port_reg_data_mux_1_nl = MUX_v_28_2_2(act_port_reg_data_59_32_sva, (PECore_RunScale_if_for_4_mul_1_cmp_4_z[38:11]),
      act_port_reg_data_and_16_cse);
  assign act_port_reg_data_mux_nl = MUX_v_28_2_2(act_port_reg_data_27_0_sva, (PECore_RunScale_if_for_4_mul_1_cmp_2_z[38:11]),
      act_port_reg_data_and_16_cse);
  assign nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun
      = signext_256_252({act_port_reg_data_mux_7_nl , (signext_32_28(act_port_reg_data_mux_6_nl))
      , (signext_32_28(act_port_reg_data_mux_5_nl)) , (signext_32_28(act_port_reg_data_mux_4_nl))
      , (signext_32_28(act_port_reg_data_mux_3_nl)) , (signext_32_28(act_port_reg_data_mux_2_nl))
      , (signext_32_28(act_port_reg_data_mux_1_nl)) , (signext_32_28(act_port_reg_data_mux_nl))});
  wire weight_port_read_out_data_mux_4_nl;
  wire weight_port_read_out_data_mux_111_nl;
  wire weight_port_read_out_data_mux_2_nl;
  wire weight_port_read_out_data_mux_110_nl;
  wire weight_port_read_out_data_mux_nl;
  wire weight_port_read_out_data_mux_109_nl;
  wire [127:0] nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign weight_port_read_out_data_mux_111_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_26_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign weight_port_read_out_data_mux_4_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1,
      weight_port_read_out_data_mux_111_nl, fsm_output);
  assign weight_port_read_out_data_mux_110_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_25_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign weight_port_read_out_data_mux_2_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1,
      weight_port_read_out_data_mux_110_nl, fsm_output);
  assign weight_port_read_out_data_mux_109_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_24_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign weight_port_read_out_data_mux_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1,
      weight_port_read_out_data_mux_109_nl, fsm_output);
  assign nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun
      = {rva_out_reg_data_127_120_sva_dfm_4_4_7_6 , rva_out_reg_data_127_120_sva_dfm_4_4_5_0
      , rva_out_reg_data_119_112_sva_dfm_4_4_7 , rva_out_reg_data_119_112_sva_dfm_4_4_6_0
      , rva_out_reg_data_111_104_sva_dfm_4_4_7 , rva_out_reg_data_111_104_sva_dfm_4_4_6_0
      , reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd , reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd_1
      , rva_out_reg_data_95_88_sva_dfm_4_4 , reg_rva_out_reg_data_87_80_sva_dfm_4_4_ftd
      , reg_rva_out_reg_data_87_80_sva_dfm_4_4_ftd_1 , rva_out_reg_data_79_72_sva_dfm_4_4
      , rva_out_reg_data_71_64_sva_dfm_4_4 , rva_out_reg_data_63_sva_dfm_4_4 , rva_out_reg_data_62_56_sva_dfm_4_4
      , rva_out_reg_data_55_48_sva_dfm_4_4 , rva_out_reg_data_47_sva_dfm_4_4 , rva_out_reg_data_46_40_sva_dfm_4_4
      , rva_out_reg_data_39_36_sva_dfm_4_4 , rva_out_reg_data_35_32_sva_dfm_4_4 ,
      PECore_PushAxiRsp_if_mux1h_17 , PECore_PushAxiRsp_if_mux1h_16 , PECore_PushAxiRsp_if_mux1h_15
      , PECore_PushAxiRsp_if_mux1h_14_6 , PECore_PushAxiRsp_if_mux1h_14_5_0 , weight_port_read_out_data_mux_4_nl
      , PECore_PushAxiRsp_if_mux1h_12_6_3 , PECore_PushAxiRsp_if_mux1h_12_2_0 , weight_port_read_out_data_mux_2_nl
      , PECore_PushAxiRsp_if_mux1h_10_6_3 , PECore_PushAxiRsp_if_mux1h_10_2_0 , weight_port_read_out_data_mux_nl};
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd31),
  .signd_b(32'sd1),
  .width_z(32'sd39),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_4_mul_1_cmp (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_4_mul_1_cmp_b[30:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_4_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_4_mul_1_cmp_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd31),
  .signd_b(32'sd1),
  .width_z(32'sd39),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_4_mul_1_cmp_1 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_4_mul_1_cmp_1_b[30:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_4_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_4_mul_1_cmp_1_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd31),
  .signd_b(32'sd1),
  .width_z(32'sd39),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_4_mul_1_cmp_2 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_4_mul_1_cmp_2_b[30:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_4_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_4_mul_1_cmp_2_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd31),
  .signd_b(32'sd1),
  .width_z(32'sd39),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_4_mul_1_cmp_3 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_4_mul_1_cmp_3_b[30:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_4_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_4_mul_1_cmp_3_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd31),
  .signd_b(32'sd1),
  .width_z(32'sd39),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_4_mul_1_cmp_4 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_4_mul_1_cmp_4_b[30:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_4_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_4_mul_1_cmp_4_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd31),
  .signd_b(32'sd1),
  .width_z(32'sd39),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_4_mul_1_cmp_5 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_4_mul_1_cmp_5_b[30:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_4_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_4_mul_1_cmp_5_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd31),
  .signd_b(32'sd1),
  .width_z(32'sd39),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_4_mul_1_cmp_6 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_4_mul_1_cmp_6_b[30:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_4_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_4_mul_1_cmp_6_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd31),
  .signd_b(32'sd1),
  .width_z(32'sd39),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_4_mul_1_cmp_7 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_4_mul_1_cmp_7_b[30:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_4_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_4_mul_1_cmp_7_z)
    );
  PECore_mgc_muladd1 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_cst(32'sd1),
  .signd_cst(32'sd0),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd11),
  .add_axb(32'sd1),
  .add_c(32'sd1),
  .add_d(32'sd1),
  .use_const(32'sd1)) PEManager_15U_GetWeightAddr_else_acc_4_cmp (
      .a(pe_config_output_counter_sva),
      .b(pe_manager_num_input_sva),
      .c(pe_config_input_counter_sva),
      .cst(1'b0),
      .z(PEManager_15U_GetWeightAddr_else_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_for_1_lshift_rg (
      .a(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a),
      .s(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_write_arbxbar_xbar_for_lshift_rg (
      .a(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a),
      .s(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s[2:0]),
      .z(weight_mem_write_arbxbar_xbar_for_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi PECore_PECoreRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(fsm_output)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi PECore_PECoreRun_input_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_oswt_pff(and_547_rmff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi PECore_PECoreRun_act_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(reg_act_port_Push_mioi_iswt0_cse),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun[255:0]),
      .act_port_Push_mioi_oswt_pff(and_549_cse)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi PECore_PECoreRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_oswt_pff(and_547_rmff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi PECore_PECoreRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun[127:0]),
      .rva_out_Push_mioi_oswt_pff(and_545_cse)
    );
  PECore_PECore_PECoreRun_wait_dp PECore_PECoreRun_wait_dp_inst (
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .ProductSum_for_acc_20_cmp_en(ProductSum_for_acc_20_cmp_en),
      .ProductSum_for_acc_19_cmp_en(ProductSum_for_acc_19_cmp_en),
      .PECoreRun_wen(PECoreRun_wen),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg(and_543_rmff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg(and_540_rmff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg(and_537_rmff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg(and_534_rmff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg(and_531_rmff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg(and_527_rmff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg(and_523_rmff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg(and_520_rmff),
      .PECore_RunScale_if_for_4_mul_1_cmp_cgo(reg_PECore_RunScale_if_for_4_mul_1_cmp_cgo_ir_7_cse),
      .PECore_RunScale_if_for_4_mul_1_cmp_cgo_ir_unreg(and_516_rmff),
      .PECore_RunScale_if_for_4_mul_1_cmp_en(PECore_RunScale_if_for_4_mul_1_cmp_en),
      .ProductSum_for_acc_20_cmp_cgo(reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_cgo_ir_cse),
      .ProductSum_for_acc_20_cmp_cgo_ir_unreg(and_514_rmff),
      .ProductSum_for_acc_19_cmp_cgo(reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_cgo_ir_cse),
      .ProductSum_for_acc_19_cmp_cgo_ir_unreg(and_511_rmff)
    );
  PECore_PECore_PECoreRun_staller PECore_PECoreRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp)
    );
  PECore_PECore_PECoreRun_PECoreRun_fsm PECore_PECoreRun_PECoreRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .fsm_output(fsm_output)
    );
  assign weight_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_88);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign weight_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_88);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign weight_mem_banks_read_1_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_90);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign weight_mem_banks_read_1_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_90);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign weight_mem_banks_read_1_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_92);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 );
  assign weight_mem_banks_read_1_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_92);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign weight_mem_banks_read_1_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_94);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 );
  assign weight_mem_banks_read_1_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_94);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign weight_mem_banks_read_1_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_96);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 );
  assign weight_mem_banks_read_1_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_96);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign weight_mem_banks_read_1_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_98);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 );
  assign weight_mem_banks_read_1_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_98);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign weight_mem_banks_read_1_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_84);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 );
  assign weight_mem_banks_read_1_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_84);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign weight_mem_banks_read_1_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_86);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 );
  assign weight_mem_banks_read_1_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_86);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign weight_mem_banks_write_if_for_if_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_171);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 );
  assign weight_mem_banks_write_if_for_if_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_171);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign weight_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_174);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 );
  assign weight_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_174);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign weight_mem_banks_write_if_for_if_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_175);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 );
  assign weight_mem_banks_write_if_for_if_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_175);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1
      = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1
      = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign weight_mem_banks_read_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_177);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 );
  assign weight_mem_banks_read_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_177);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign weight_mem_banks_write_if_for_if_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_178);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 );
  assign weight_mem_banks_write_if_for_if_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_178);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2
      = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2
      = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign weight_mem_banks_read_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_181);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 );
  assign weight_mem_banks_read_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_181);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign weight_mem_banks_write_if_for_if_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_182);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 );
  assign weight_mem_banks_write_if_for_if_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_182);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3
      = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3
      = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign weight_mem_banks_read_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_185);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 );
  assign weight_mem_banks_read_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_185);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign weight_mem_banks_write_if_for_if_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_187);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 );
  assign weight_mem_banks_write_if_for_if_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_187);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4
      = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4
      = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign weight_mem_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_190);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 );
  assign weight_mem_banks_read_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_190);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign weight_mem_banks_write_if_for_if_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_191);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 );
  assign weight_mem_banks_write_if_for_if_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_191);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5
      = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5
      = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign weight_mem_banks_read_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_194);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 );
  assign weight_mem_banks_read_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_194);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign weight_mem_banks_write_if_for_if_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_196);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 );
  assign weight_mem_banks_write_if_for_if_mux_33_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_196);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6
      = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6
      = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign weight_mem_banks_read_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_198);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 );
  assign weight_mem_banks_read_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_198);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign weight_mem_banks_write_if_for_if_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_200);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 );
  assign weight_mem_banks_write_if_for_if_mux_37_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_200);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7
      = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7
      = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign weight_mem_banks_read_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_202);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 );
  assign weight_mem_banks_read_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_202);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign input_mem_banks_write_1_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_212);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 );
  assign input_mem_banks_write_1_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_212);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8
      = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_3 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8
      = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign input_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_209);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 );
  assign input_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_209);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign input_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_219);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 );
  assign input_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_219);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9
      = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_1 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9
      = input_mem_banks_write_if_for_if_mux_1_cse;
  assign input_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_222);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 );
  assign input_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_222);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign and_511_rmff = (and_dcpl_507 | ((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_7 & while_stage_0_9)) & fsm_output;
  assign and_514_rmff = (and_dcpl_35 | and_dcpl_507) & fsm_output;
  assign and_516_rmff = (~(((~ while_stage_0_9) | PECore_RunMac_PECore_RunMac_if_and_svs_st_7
      | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8)
      | (~ while_stage_0_10) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)))
      & fsm_output;
  assign or_359_nl = weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | and_tmp_4;
  assign or_358_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3)))
      | and_tmp_4;
  assign mux_100_nl = MUX_s_1_2_2(or_359_nl, or_358_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_101_nl = MUX_s_1_2_2(and_tmp_4, mux_100_nl, while_stage_0_7);
  assign and_520_rmff = (mux_101_nl | and_dcpl_514) & fsm_output;
  assign or_363_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | and_tmp_5;
  assign or_362_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3)))
      | and_tmp_5;
  assign mux_103_nl = MUX_s_1_2_2(or_363_nl, or_362_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_104_nl = MUX_s_1_2_2(and_tmp_5, mux_103_nl, while_stage_0_7);
  assign and_523_rmff = (mux_104_nl | and_dcpl_516) & fsm_output;
  assign or_370_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_6;
  assign or_369_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2)))
      | and_tmp_6;
  assign mux_106_nl = MUX_s_1_2_2(or_370_nl, or_369_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_107_nl = MUX_s_1_2_2(and_tmp_6, mux_106_nl, while_stage_0_6);
  assign and_527_rmff = (mux_107_nl | and_dcpl_191) & fsm_output;
  assign or_376_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_7;
  assign or_836_nl = (~((~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1)) | and_tmp_7;
  assign mux_109_nl = MUX_s_1_2_2(or_376_nl, or_836_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_110_nl = MUX_s_1_2_2(and_tmp_7, mux_109_nl, while_stage_0_6);
  assign and_531_rmff = (mux_110_nl | and_dcpl_187) & fsm_output;
  assign or_382_nl = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_8;
  assign or_837_nl = (~((~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1)) | and_tmp_8;
  assign mux_113_nl = MUX_s_1_2_2(or_382_nl, or_837_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_114_nl = MUX_s_1_2_2(and_tmp_8, mux_113_nl, while_stage_0_6);
  assign and_534_rmff = (mux_114_nl | and_dcpl_182) & fsm_output;
  assign or_388_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_9;
  assign or_838_nl = (~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1)) | and_tmp_9;
  assign mux_116_nl = MUX_s_1_2_2(or_388_nl, or_838_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_117_nl = MUX_s_1_2_2(and_tmp_9, mux_116_nl, while_stage_0_6);
  assign and_537_rmff = (mux_117_nl | and_dcpl_178) & fsm_output;
  assign or_394_nl = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_10;
  assign or_839_nl = (~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1)) | and_tmp_10;
  assign mux_119_nl = MUX_s_1_2_2(or_394_nl, or_839_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_120_nl = MUX_s_1_2_2(and_tmp_10, mux_119_nl, while_stage_0_6);
  assign and_540_rmff = (mux_120_nl | and_dcpl_175) & fsm_output;
  assign or_400_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_11;
  assign or_399_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse)))
      | and_tmp_11;
  assign mux_123_nl = MUX_s_1_2_2(or_400_nl, or_399_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_124_nl = MUX_s_1_2_2(and_tmp_11, mux_123_nl, while_stage_0_6);
  assign and_543_rmff = (mux_124_nl | and_dcpl_171) & fsm_output;
  assign and_1075_nl = PECore_UpdateFSM_switch_lp_nor_7_itm_1 & PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      & pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign and_755_nl = pe_config_is_zero_first_sva & PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      & pe_manager_zero_active_sva;
  assign mux_433_itm = MUX_s_1_2_2(and_1075_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_755_nl);
  assign and_759_nl = start_PopNB_mioi_data_rsc_z_mxwt & start_PopNB_mioi_return_rsc_z_mxwt
      & PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign mux_133_nl = MUX_s_1_2_2(mux_433_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_759_nl);
  assign mux_129_nl = MUX_s_1_2_2(mux_433_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_754_cse);
  assign mux_134_nl = MUX_s_1_2_2(mux_133_nl, mux_129_nl, or_407_cse);
  assign mux_428_nl = MUX_s_1_2_2(mux_433_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_754_cse);
  assign or_405_nl = pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]);
  assign mux_130_nl = MUX_s_1_2_2(mux_428_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_405_nl);
  assign or_404_nl = (state_2_1_sva!=2'b10) | state_0_sva;
  assign mux_131_nl = MUX_s_1_2_2(mux_130_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_404_nl);
  assign mux_132_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_nor_7_itm_1, mux_131_nl,
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign mux_135_nl = MUX_s_1_2_2(mux_134_nl, mux_132_nl, PECore_UpdateFSM_switch_lp_equal_tmp_5_1);
  assign mux_136_cse = MUX_s_1_2_2(mux_135_nl, state_0_sva, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_137_nl = MUX_s_1_2_2(or_407_cse, mux_136_cse, while_stage_0_3);
  assign or_403_nl = while_stage_0_3 | (state_2_1_sva!=2'b00) | state_0_sva;
  assign or_402_nl = (state_2_1_sva_dfm_1!=2'b00);
  assign mux_138_nl = MUX_s_1_2_2(mux_137_nl, or_403_nl, or_402_nl);
  assign and_547_rmff = (~ mux_138_nl) & and_dcpl_213;
  assign PECore_DecodeAxiRead_switch_lp_and_2_cse = PECoreRun_wen & and_dcpl_8;
  assign rva_out_reg_data_and_23_cse = PECoreRun_wen & and_dcpl_8 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_8) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8)
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 | rva_in_reg_rw_sva_st_8));
  assign rva_out_reg_data_and_128_enex5 = rva_out_reg_data_and_23_cse & reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  assign rva_out_reg_data_and_129_enex5 = rva_out_reg_data_and_23_cse & reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_130_enex5 = rva_out_reg_data_and_23_cse & reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_26_cse = PECoreRun_wen & and_dcpl_7;
  assign rva_out_reg_data_and_131_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_132_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_133_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_95_88_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_134_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_135_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_136_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_79_72_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_137_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_71_64_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_138_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_139_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_140_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_141_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_142_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo;
  assign input_mem_banks_read_read_data_and_cse = PECoreRun_wen & and_dcpl_7 & (~
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6) & input_read_req_valid_lpi_1_dfm_1_8;
  assign weight_port_read_out_data_and_122_cse = PECoreRun_wen & and_dcpl_6 & (~
      rva_in_reg_rw_sva_st_1_8) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  assign rva_out_reg_data_and_cse = PECoreRun_wen & (~((~(while_stage_0_11 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9))
      | rva_in_reg_rw_sva_9 | (~ fsm_output)));
  assign input_mem_banks_read_read_data_and_35_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo;
  assign weight_port_read_out_data_and_213_enex5 = weight_port_read_out_data_and_122_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_3_enexo;
  assign input_mem_banks_read_read_data_and_36_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_37_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_38_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo;
  assign rva_in_reg_rw_and_cse = PECoreRun_wen & while_stage_0_10;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_cse = PECoreRun_wen & and_dcpl_6
      & (~(rva_in_reg_rw_sva_st_1_8 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6))
      & (~(rva_in_reg_rw_sva_8 | input_read_req_valid_lpi_1_dfm_1_8)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  assign PECore_PushOutput_if_and_cse = PECoreRun_wen & and_dcpl_24;
  assign or_851_nl = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_8) | PECore_RunMac_PECore_RunMac_if_and_svs_8
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  assign mux_436_nl = MUX_s_1_2_2(not_tmp_488, or_tmp_484, or_851_nl);
  assign mux_435_nl = MUX_s_1_2_2(not_tmp_488, or_tmp_484, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nor_nl = ~(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8));
  assign mux_437_nl = MUX_s_1_2_2(mux_436_nl, mux_435_nl, nor_nl);
  assign and_1086_cse = mux_437_nl & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)
      & while_stage_0_11 & PECoreRun_wen;
  assign PECore_RunScale_if_and_cse = PECoreRun_wen & and_dcpl_24 & (PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8
      | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8));
  assign accum_vector_data_and_cse = rva_in_reg_rw_and_cse & while_stage_0_10;
  assign rva_in_reg_rw_and_2_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & while_stage_0_9;
  assign and_1125_cse = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | accum_vector_operator_1_for_asn_115_itm_7);
  assign and_1140_cse = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | accum_vector_operator_1_for_asn_100_itm_7);
  assign and_1155_cse = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | accum_vector_operator_1_for_asn_85_itm_7);
  assign and_1170_cse = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | accum_vector_operator_1_for_asn_73_itm_7);
  assign and_1188_cse = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | accum_vector_operator_1_for_asn_55_itm_7);
  assign and_1203_cse = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | accum_vector_operator_1_for_asn_43_itm_7);
  assign and_1221_cse = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | accum_vector_operator_1_for_asn_25_itm_7);
  assign and_1236_cse = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | accum_vector_operator_1_for_asn_10_itm_7);
  assign accum_vector_operator_1_for_and_cse = PECoreRun_wen & and_dcpl_29;
  assign while_if_and_6_cse = PECoreRun_wen & while_stage_0_9;
  assign PECore_RunMac_if_and_2_cse = PECoreRun_wen & and_dcpl_33;
  assign while_if_and_7_cse = PECoreRun_wen & while_stage_0_8;
  assign ProductSum_for_and_cse = PECoreRun_wen & and_dcpl_35;
  assign input_mem_banks_read_1_read_data_and_enex5 = ProductSum_for_and_cse & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  assign weight_port_read_out_data_7_0_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]),
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9, weight_port_read_out_data_7_0_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_100_itm_1 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_3_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]), weight_port_read_out_data_7_3_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_100_itm_1 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_2_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]), weight_port_read_out_data_7_2_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_100_itm_1 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_5_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]), weight_port_read_out_data_7_5_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_4_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]), weight_port_read_out_data_7_4_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_7_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]), weight_port_read_out_data_7_7_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_6_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]), weight_port_read_out_data_7_6_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_9_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]), weight_port_read_out_data_7_9_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_8_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]), weight_port_read_out_data_7_8_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_11_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]), weight_port_read_out_data_7_11_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_10_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]), weight_port_read_out_data_7_10_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_100_itm_1 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_13_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), weight_port_read_out_data_7_13_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_12_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]), weight_port_read_out_data_7_12_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_15_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), weight_port_read_out_data_7_15_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_14_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), weight_port_read_out_data_7_14_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_15_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), weight_port_read_out_data_5_15_sva_dfm_1_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , weight_mem_run_3_for_5_and_12_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_weight_mem_run_3_for_5_and_14_itm_1_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , reg_weight_mem_run_3_for_5_and_16_itm_1_cse , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_14_sva_dfm_1_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), weight_port_read_out_data_5_14_sva_dfm_1_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , weight_mem_run_3_for_5_and_7_itm_1 , reg_weight_mem_run_3_for_5_and_16_itm_1_cse
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_and_cse = PECoreRun_wen & (~(or_dcpl_243 | (~
      weight_mem_run_3_for_land_5_lpi_1_dfm_3)));
  assign weight_port_read_out_data_and_214_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  assign data_in_tmp_operator_2_for_and_cse = PECoreRun_wen & weight_mem_run_3_for_land_5_lpi_1_dfm_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7;
  assign weight_mem_run_3_for_aelse_and_cse = PECoreRun_wen & while_stage_0_7;
  assign weight_port_read_out_data_and_215_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001;
  assign weight_port_read_out_data_and_216_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002;
  assign weight_port_read_out_data_and_217_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003;
  assign weight_port_read_out_data_and_218_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004;
  assign weight_port_read_out_data_and_219_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005;
  assign weight_port_read_out_data_and_220_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006;
  assign weight_port_read_out_data_and_221_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007;
  assign weight_port_read_out_data_and_222_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008;
  assign weight_port_read_out_data_and_223_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009;
  assign weight_port_read_out_data_and_224_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010;
  assign weight_port_read_out_data_and_225_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011;
  assign weight_port_read_out_data_and_226_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012;
  assign weight_port_read_out_data_and_227_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013;
  assign weight_port_read_out_data_and_228_enex5 = weight_port_read_out_data_and_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014;
  assign weight_port_read_out_data_and_15_enex5 = PECoreRun_wen & (~(or_dcpl_243
      | (~ weight_mem_run_3_for_land_4_lpi_1_dfm_3) | (~ fsm_output))) & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7) | (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)) & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  assign weight_port_read_out_data_and_16_cse = PECoreRun_wen & (~(or_dcpl_243 |
      (~ weight_mem_run_3_for_land_3_lpi_1_dfm_3)));
  assign weight_port_read_out_data_and_229_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  assign data_in_tmp_operator_2_for_and_16_cse = PECoreRun_wen & weight_mem_run_3_for_land_3_lpi_1_dfm_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7;
  assign weight_port_read_out_data_and_230_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001;
  assign weight_port_read_out_data_and_231_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002;
  assign weight_port_read_out_data_and_232_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003;
  assign weight_port_read_out_data_and_233_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004;
  assign weight_port_read_out_data_and_234_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005;
  assign weight_port_read_out_data_and_235_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006;
  assign weight_port_read_out_data_and_236_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007;
  assign weight_port_read_out_data_and_237_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008;
  assign weight_port_read_out_data_and_238_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009;
  assign weight_port_read_out_data_and_239_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010;
  assign weight_port_read_out_data_and_240_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011;
  assign weight_port_read_out_data_and_241_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012;
  assign weight_port_read_out_data_and_242_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013;
  assign weight_port_read_out_data_and_243_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014;
  assign weight_port_read_out_data_and_31_enex5 = PECoreRun_wen & (~(or_dcpl_243
      | (~ weight_mem_run_3_for_land_2_lpi_1_dfm_3))) & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  assign weight_mem_run_3_for_5_and_159_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_161_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_cse = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_173_cse = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_174_cse = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_176_cse = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_178_cse = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_179_cse = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign or_931_cse = (~ weight_mem_run_3_for_land_1_lpi_1_dfm_2) | (~ while_stage_0_6)
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  assign or_928_cse = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)
      | (~ while_stage_0_6) | PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  assign PECore_RunMac_if_and_3_cse = PECoreRun_wen & and_dcpl_40;
  assign and_572_cse = nor_tmp_2 & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2:1]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      | (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1:0]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_or_2_cse = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3) | ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_1006_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_dcpl);
  assign and_1007_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_2_cse & (~
      or_dcpl);
  assign and_1008_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      & (~ or_dcpl);
  assign and_1009_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      & (~ or_dcpl);
  assign and_1010_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      & (~ or_dcpl);
  assign and_1011_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      & (~ or_dcpl);
  assign nor_506_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl);
  assign rva_in_reg_rw_and_3_cse = PECoreRun_wen & and_dcpl_54;
  assign weight_mem_banks_read_1_read_data_and_8_cse = PECoreRun_wen & and_dcpl_55;
  assign ProductSum_for_and_8_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign input_mem_banks_read_1_read_data_and_5_enex5 = ProductSum_for_and_8_cse
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  assign weight_mem_run_3_for_aelse_and_4_cse = PECoreRun_wen & while_stage_0_6;
  assign weight_port_read_out_data_and_137_cse = PECoreRun_wen & (~(or_dcpl_252 |
      (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2) | (~ fsm_output))) & (or_dcpl_12
      | (~ weight_mem_run_3_for_land_4_lpi_1_dfm_1));
  assign xor_1_cse = (weight_read_addrs_7_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[2]);
  assign and_1279_cse = (xor_1_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign or_939_cse = and_1279_cse | weight_mem_run_3_for_5_and_31_itm_2 | weight_mem_run_3_for_5_and_30_itm_2
      | weight_mem_run_3_for_5_and_28_itm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse = PECoreRun_wen
      & and_dcpl_55 & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_375_cse = PECoreRun_wen
      & and_dcpl_55 & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_379_cse = PECoreRun_wen
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_4_lpi_1_dfm_1) & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_380_cse = PECoreRun_wen
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1 & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_382_cse = PECoreRun_wen
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_2_lpi_1_dfm_1) & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_cse = PECoreRun_wen
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_2 & while_stage_0_6;
  assign weight_read_addrs_and_5_cse = PECoreRun_wen & (((~ ProductSum_for_asn_69_itm_3)
      & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1)
      | (weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
      & (~ ProductSum_for_asn_56_itm_3))) & and_dcpl_76;
  assign weight_read_addrs_and_28_enex5 = weight_read_addrs_and_5_cse & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_2_cse = PECoreRun_wen & and_dcpl_84;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_2_cse
      & (reg_weight_read_addrs_3_lpi_1_dfm_1_enexo | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3_enexo
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo);
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_4_cse = PECoreRun_wen & and_dcpl_86;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_4_cse
      & (reg_weight_read_addrs_3_lpi_1_dfm_1_enexo_1 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1
      | reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo);
  assign while_if_and_10_cse = PECoreRun_wen & while_stage_0_5;
  assign weight_mem_read_arbxbar_arbiters_next_and_cse = PECoreRun_wen & fsm_output;
  assign weight_mem_read_arbxbar_arbiters_next_and_48_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_107_cse | or_237_cse);
  assign weight_mem_read_arbxbar_arbiters_next_and_54_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_114_cse | or_237_cse);
  assign weight_mem_read_arbxbar_arbiters_next_and_60_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_121_cse | or_237_cse);
  assign weight_mem_read_arbxbar_arbiters_next_and_66_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((nor_294_cse & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) |
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]))) & nor_297_cse) | or_237_cse);
  assign weight_mem_read_arbxbar_arbiters_next_and_72_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_135_cse | or_237_cse);
  assign weight_mem_read_arbxbar_arbiters_next_and_78_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_142_cse | or_237_cse);
  assign weight_mem_read_arbxbar_arbiters_next_and_84_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((nor_306_cse & nor_307_cse & nor_308_cse & nor_309_cse) | or_237_cse);
  assign weight_mem_read_arbxbar_arbiters_next_and_90_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_156_cse | or_237_cse);
  assign weight_read_addrs_and_7_cse = PECoreRun_wen & while_stage_0_4;
  assign weight_write_data_data_and_cse = PECoreRun_wen & ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7:6]!=2'b00))
      & and_dcpl_155;
  assign weight_write_data_data_and_48_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_49_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_50_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_51_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_52_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_53_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_54_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_55_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_56_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_57_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_58_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_59_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_60_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_61_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_62_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_63_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_addrs_and_enex5 = weight_write_data_data_and_cse & reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
      = PECoreRun_wen & and_dcpl_162;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 & and_dcpl_162;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 & and_dcpl_162;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12 & and_dcpl_162;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_25_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13 & and_dcpl_162;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14 & and_dcpl_162;
  assign Arbiter_8U_Roundrobin_pick_1_and_15_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8
      & and_dcpl_162;
  assign weight_mem_read_arbxbar_xbar_requests_transpose_and_13_cse = PECoreRun_wen
      & and_dcpl_155;
  assign Arbiter_8U_Roundrobin_pick_and_cse = PECoreRun_wen & (while_stage_0_4 |
      and_dcpl_576) & fsm_output & or_237_cse;
  assign Arbiter_8U_Roundrobin_pick_1_and_22_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9
      & and_dcpl_162;
  assign Arbiter_8U_Roundrobin_pick_1_and_64_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15
      & and_dcpl_162;
  assign weight_write_data_data_and_16_cse = PECoreRun_wen & and_dcpl_205;
  assign weight_write_data_data_and_64_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_65_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_66_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_67_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_68_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_69_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_70_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_71_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_72_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_73_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_74_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_75_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_76_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_77_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_78_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_79_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  assign weight_write_addrs_and_2_enex5 = weight_write_data_data_and_16_cse & reg_pe_manager_base_input_enexo;
  assign PECore_DecodeAxiWrite_switch_lp_and_2_cse = PECoreRun_wen & while_stage_0_3;
  assign weight_read_addrs_and_29_enex5 = weight_write_data_data_and_16_cse & reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  assign state_and_cse = weight_mem_read_arbxbar_arbiters_next_and_cse & nand_91_cse;
  assign and_1287_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & while_stage_0_3;
  assign pe_config_num_manager_and_cse = PECoreRun_wen & (~(or_dcpl_271 | or_dcpl_270
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]))));
  assign rva_in_reg_rw_and_5_cse = PECoreRun_wen & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign PECore_UpdateFSM_switch_lp_and_9_cse = PECoreRun_wen & and_dcpl_213;
  assign or_945_cse = (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign nor_571_cse = ~((~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1);
  assign and_1600_cse = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  assign pe_config_UpdateManagerCounter_if_if_and_enex5 = PECoreRun_wen & reg_pe_config_num_output_enexo;
  assign PECore_DecodeAxiRead_switch_lp_and_cse = PECoreRun_wen & (~(nand_91_cse
      | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
  assign PECore_DecodeAxiWrite_switch_lp_and_cse = PECoreRun_wen & (~ or_dcpl_270);
  assign weight_port_read_out_data_and_138_cse = PECoreRun_wen & and_dcpl_224 & while_stage_0_9
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  assign weight_port_read_out_data_and_244_enex5 = weight_port_read_out_data_and_138_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_2_enexo;
  assign weight_port_read_out_data_and_245_enex5 = weight_port_read_out_data_and_138_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  assign weight_port_read_out_data_and_246_enex5 = weight_port_read_out_data_and_138_cse
      & reg_weight_port_read_out_data_0_2_sva_dfm_2_1_enexo;
  assign and_1023_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_2_cse & (~
      or_dcpl_329);
  assign and_1024_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      & (~ or_dcpl_329);
  assign and_1025_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      & (~ or_dcpl_329);
  assign and_1026_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1
      & (~ or_dcpl_329);
  assign and_1027_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      & (~ or_dcpl_329);
  assign nor_508_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl_329);
  assign weight_mem_banks_load_store_for_else_and_1_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_mem_banks_load_store_for_else_and_2_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_read_addrs_and_17_cse = PECoreRun_wen & weight_mem_run_3_for_land_3_lpi_1_dfm_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign weight_port_read_out_data_and_143_cse = PECoreRun_wen & (~(or_dcpl_251 |
      (~ fsm_output))) & (or_dcpl_12 | (~ weight_mem_run_3_for_land_7_lpi_1_dfm_1));
  assign weight_port_read_out_data_and_158_cse = PECoreRun_wen & (~(or_dcpl_253 |
      (~ fsm_output))) & (or_dcpl_12 | (~ weight_mem_run_3_for_land_6_lpi_1_dfm_1_1));
  assign weight_port_read_out_data_and_185_cse = PECoreRun_wen & (~(or_dcpl_255 |
      (~ fsm_output))) & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_run_3_for_land_2_lpi_1_dfm_1) | (~ while_stage_0_6));
  assign weight_port_read_out_data_and_199_cse = PECoreRun_wen & (while_and_1243_cse
      | while_and_40_tmp) & while_stage_0_7 & fsm_output & (~(mux_15_itm & while_stage_0_6));
  assign nor_573_cse = ~((weight_read_addrs_7_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_467_nl = MUX_s_1_2_2((weight_read_addrs_7_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_7_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_7_lpi_1_dfm_3_2_0[0]);
  assign mux_468_cse = MUX_s_1_2_2(mux_467_nl, nor_573_cse, weight_read_addrs_7_lpi_1_dfm_3_2_0[2]);
  assign and_1327_cse = (mux_468_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign and_1332_cse = (xor_1_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign and_1352_cse = (mux_468_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign and_1363_cse = (and_1327_cse | or_dcpl_408 | or_dcpl_394) & and_dcpl_958
      & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign nor_582_cse = ~((weight_read_addrs_5_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_485_nl = MUX_s_1_2_2((weight_read_addrs_5_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_5_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_5_lpi_1_dfm_3_2_0[0]);
  assign mux_486_nl = MUX_s_1_2_2(mux_485_nl, nor_582_cse, weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign and_1397_cse = (mux_486_nl | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_384_cse = PECoreRun_wen
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_6_lpi_1_dfm_1_1) & while_stage_0_6;
  assign nor_352_cse = ~(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign weight_read_addrs_and_19_cse = PECoreRun_wen & and_dcpl_82;
  assign weight_read_addrs_and_20_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse
      & and_dcpl_248;
  assign or_222_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]);
  assign and_743_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_4_sva;
  assign and_742_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_3_sva;
  assign and_744_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  assign mux_592_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp,
      mux_tmp_42, and_743_cse);
  assign mux_47_itm = MUX_s_1_2_2(mux_tmp_42, mux_592_nl, and_742_cse);
  assign and_745_cse = (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 |
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign or_237_cse = (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_30_cse
      = weight_mem_read_arbxbar_arbiters_next_and_cse & or_237_cse;
  assign operator_15_false_1_and_cse = PECoreRun_wen & (~(and_107_cse | or_237_cse));
  assign PEManager_15U_PEManagerWrite_and_enex5 = PECoreRun_wen & reg_rva_in_reg_rw_sva_st_1_1_cse
      & (~ PECore_DecodeAxiWrite_switch_lp_equal_tmp_1) & (~ PECore_DecodeAxiWrite_switch_lp_nor_tmp_1)
      & PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 & (~ PECore_DecodeAxiWrite_switch_lp_equal_tmp_2)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_in_reg_data_sva_1_enexo;
  assign pe_manager_num_input_and_cse = PECoreRun_wen & (~(or_dcpl_271 | nand_91_cse
      | or_dcpl_305));
  assign pe_config_is_valid_and_cse = PECoreRun_wen & (~(PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1
      | PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (~ nand_91_cse);
  assign nor_589_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:10]!=2'b00));
  assign nor_524_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])));
  assign while_if_and_14_cse = PECoreRun_wen & and_cse;
  assign rva_in_reg_rw_and_6_cse = PECoreRun_wen & and_dcpl_76;
  assign rva_in_reg_rw_and_7_cse = PECoreRun_wen & and_dcpl_262;
  assign ProductSum_for_and_14_cse = PECoreRun_wen & PECore_RunMac_PECore_RunMac_if_and_svs_st_3
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_404_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_408_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_152_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign input_mem_banks_read_read_data_and_9_cse = PECoreRun_wen & and_dcpl_277
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5) & input_read_req_valid_lpi_1_dfm_1_7;
  assign input_mem_banks_read_read_data_and_39_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_40_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_41_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_42_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse = PECoreRun_wen & and_dcpl_224
      & (~ rva_in_reg_rw_sva_7) & while_stage_0_9 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5) & (~ input_read_req_valid_lpi_1_dfm_1_7);
  assign input_mem_banks_read_1_read_data_and_6_enex5 = ProductSum_for_and_14_cse
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  assign or_260_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
      | and_747_cse | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp
      | and_749_cse;
  assign weight_read_addrs_and_30_enex5 = weight_write_data_data_and_16_cse & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  assign input_read_req_valid_and_1_cse = PECoreRun_wen & and_dcpl_277;
  assign PECore_DecodeAxiRead_switch_lp_and_7_cse = PECoreRun_wen & and_dcpl_290
      & while_stage_0_9 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5)
      & (~ input_read_req_valid_lpi_1_dfm_1_7);
  assign rva_out_reg_data_and_41_cse = PECoreRun_wen & and_dcpl_290 & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_7
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7))
      & (~ rva_in_reg_rw_sva_st_7) & while_stage_0_9 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6
      & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 | input_read_req_valid_lpi_1_dfm_1_7));
  assign rva_out_reg_data_and_143_enex5 = rva_out_reg_data_and_41_cse & reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_144_enex5 = rva_out_reg_data_and_41_cse & reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_145_enex5 = rva_out_reg_data_and_41_cse & reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  assign weight_port_read_out_data_and_247_enex5 = weight_port_read_out_data_and_138_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_2_1_enexo;
  assign rva_out_reg_data_and_146_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_147_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_148_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_149_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_150_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_151_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_127_120_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_152_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_119_112_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_153_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_111_104_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_154_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_95_88_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_155_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_79_72_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_156_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_71_64_sva_dfm_4_2_enexo;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_235_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[127:120]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_235_nl);
  assign weight_mem_banks_load_store_for_else_and_4_cse = PECoreRun_wen & while_stage_0_6
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_236_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[119:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_236_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_237_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[111:104]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_237_nl);
  assign weight_mem_banks_load_store_for_else_and_56_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 & and_dcpl_54;
  assign and_1030_cse = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])
      & (~ or_dcpl_333);
  assign and_1031_cse = and_dcpl_637 & (~ or_dcpl_333);
  assign and_1032_cse = and_dcpl_638 & (~ or_dcpl_333);
  assign mux_66_nl = MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]),
      (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2])), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign nor_320_nl = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])
      | (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]));
  assign mux_67_nl = MUX_s_1_2_2(mux_66_nl, nor_320_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign weight_mem_banks_load_store_for_else_and_57_cse = PECoreRun_wen & mux_67_nl
      & and_572_cse;
  assign weight_mem_banks_load_store_for_else_and_62_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_mem_banks_load_store_for_else_and_64_cse = PECoreRun_wen & and_572_cse
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_1;
  assign weight_mem_banks_load_store_for_else_and_67_cse = PECoreRun_wen & and_dcpl_54
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_1;
  assign weight_mem_write_arbxbar_xbar_for_empty_and_enex5 = rva_in_reg_rw_and_6_cse
      & reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  assign and_315_cse = PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]);
  assign rva_in_reg_rw_and_10_cse = PECoreRun_wen & and_dcpl_47;
  assign ProductSum_for_and_22_cse = PECoreRun_wen & or_tmp_8 & while_stage_0_4;
  assign ProductSum_for_and_26_cse = PECoreRun_wen & and_dcpl_323 & while_stage_0_4;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_410_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_6_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign pe_manager_base_weight_and_5_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse
      & and_dcpl_248;
  assign pe_manager_base_weight_and_6_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_3_or_cse
      & and_dcpl_248;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_158_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_1_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign input_mem_banks_read_read_data_and_18_cse = PECoreRun_wen & and_dcpl_353
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4) & input_read_req_valid_lpi_1_dfm_1_6;
  assign input_mem_banks_read_read_data_and_43_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_weight_mem_run_3_for_5_mux_11_itm_1_1_enexo;
  assign input_mem_banks_read_read_data_and_44_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_weight_mem_run_3_for_5_mux_107_itm_1_1_enexo;
  assign input_mem_banks_read_read_data_and_45_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_weight_mem_run_3_for_5_mux_108_itm_1_1_enexo;
  assign input_mem_banks_read_read_data_and_46_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_weight_mem_run_3_for_5_mux_109_itm_1_1_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse = PECoreRun_wen & and_dcpl_352
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 & while_stage_0_8 & and_dcpl_356;
  assign input_mem_banks_read_1_read_data_and_7_enex5 = ProductSum_for_and_26_cse
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  assign input_read_req_valid_and_2_cse = PECoreRun_wen & and_dcpl_353;
  assign PECore_DecodeAxiRead_switch_lp_and_11_cse = PECoreRun_wen & and_dcpl_353
      & and_dcpl_356;
  assign rva_out_reg_data_and_57_cse = PECoreRun_wen & and_dcpl_352 & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_6)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 & (~ rva_in_reg_rw_sva_st_6)
      & while_stage_0_8 & and_dcpl_356 & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6));
  assign rva_out_reg_data_and_157_enex5 = rva_out_reg_data_and_57_cse & reg_weight_mem_run_3_for_5_mux_12_itm_1_1_enexo;
  assign rva_out_reg_data_and_158_enex5 = rva_out_reg_data_and_57_cse & reg_weight_mem_run_3_for_5_mux_111_itm_1_1_enexo;
  assign rva_out_reg_data_and_159_enex5 = rva_out_reg_data_and_57_cse & reg_weight_mem_run_3_for_5_mux_110_itm_1_1_enexo;
  assign rva_out_reg_data_and_160_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_161_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_162_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_163_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_164_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_165_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_95_88_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_166_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_79_72_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_167_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_71_64_sva_dfm_4_1_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_3_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp;
  assign PECore_RunMac_if_and_8_cse = PECoreRun_wen & and_dcpl_206;
  assign ProductSum_for_and_30_cse = PECoreRun_wen & while_and_4_cse;
  assign input_mem_banks_read_read_data_and_27_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7 & (~(rva_in_reg_rw_sva_st_1_5 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse = PECoreRun_wen & (~ rva_in_reg_rw_sva_5)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & and_dcpl_382;
  assign input_read_req_valid_and_3_cse = PECoreRun_wen & and_dcpl_47 & (~ rva_in_reg_rw_sva_st_1_5);
  assign PECore_DecodeAxiRead_switch_lp_and_15_cse = PECoreRun_wen & (~(rva_in_reg_rw_sva_5
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & and_dcpl_382;
  assign nand_76_cse = ~(while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6);
  assign and_1442_cse = (~(((~(nand_76_cse | rva_in_reg_rw_sva_6 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)) | rva_in_reg_rw_sva_st_1_5)
      & rva_in_reg_rw_sva_5)) & weight_mem_run_3_for_aelse_and_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign nor_375_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp | (~
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp));
  assign nor_374_cse = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | ProductSum_for_asn_56_itm_1);
  assign and_1463_cse = ((~(while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5))
      | rva_in_reg_rw_sva_5) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
      & while_stage_0_8 & (~ rva_in_reg_rw_sva_6) & weight_mem_read_arbxbar_arbiters_next_and_cse;
  assign or_328_nl = rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | nand_91_cse;
  assign or_327_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign mux_87_cse = MUX_s_1_2_2(or_328_nl, or_327_nl, while_stage_0_3);
  assign mux_88_nl = MUX_s_1_2_2(mux_87_cse, or_1098_cse, while_stage_0_5);
  assign mux_89_nl = MUX_s_1_2_2(mux_88_nl, or_1097_cse, while_stage_0_6);
  assign or_326_nl = (~ while_stage_0_5) | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | rva_in_reg_rw_sva_3;
  assign mux_85_nl = MUX_s_1_2_2(or_326_nl, or_1097_cse, while_stage_0_6);
  assign mux_83_nl = MUX_s_1_2_2(reg_rva_in_reg_rw_sva_2_cse, or_1098_cse, while_stage_0_5);
  assign mux_84_nl = MUX_s_1_2_2(mux_83_nl, or_1097_cse, while_stage_0_6);
  assign mux_86_nl = MUX_s_1_2_2(mux_85_nl, mux_84_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign mux_90_nl = MUX_s_1_2_2(mux_89_nl, mux_86_nl, while_stage_0_4);
  assign rva_out_reg_data_and_93_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7 & fsm_output & mux_90_nl;
  assign nand_91_cse = ~(rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse);
  assign or_1098_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | rva_in_reg_rw_sva_3;
  assign or_1097_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | rva_in_reg_rw_sva_4;
  assign or_1099_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | reg_rva_in_reg_rw_sva_2_cse;
  assign mux_505_nl = MUX_s_1_2_2(mux_87_cse, or_1099_nl, while_stage_0_4);
  assign mux_506_nl = MUX_s_1_2_2(mux_505_nl, or_1098_cse, while_stage_0_5);
  assign mux_507_nl = MUX_s_1_2_2(mux_506_nl, or_1097_cse, while_stage_0_6);
  assign and_1488_cse = mux_507_nl & and_dcpl_958 & PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~ rva_in_reg_rw_sva_5);
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse = PECoreRun_wen & (~(rva_in_reg_rw_sva_st_1_4
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3
      & (~ rva_in_reg_rw_sva_4) & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign PECore_RunMac_if_and_10_cse = PECoreRun_wen & and_dcpl_55 & ((~ PECore_UpdateFSM_switch_lp_equal_tmp_2_4)
      | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse);
  assign mux_92_nl = MUX_s_1_2_2(or_tmp_24, and_tmp_1, weight_mem_run_3_for_land_6_lpi_1_dfm_1_1);
  assign PECore_DecodeAxiRead_switch_lp_and_19_cse = PECoreRun_wen & (~ mux_92_nl)
      & while_stage_0_6;
  assign or_511_nl = state_0_sva | (state_2_1_sva!=2'b01) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign and_682_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & (state_0_sva | (state_2_1_sva_dfm_1[1]) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign mux_167_nl = MUX_s_1_2_2(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1,
      and_682_nl, state_2_1_sva_dfm_1[0]);
  assign mux_168_nl = MUX_s_1_2_2(or_511_nl, mux_167_nl, while_stage_0_3);
  assign and_724_cse = PECoreRun_wen & (~ mux_168_nl);
  assign nor_384_cse = ~(PECore_UpdateFSM_switch_lp_equal_tmp_3_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign accum_vector_operator_1_for_and_45_cse = PECoreRun_wen & (~((~(and_dcpl_415
      & nor_329_cse)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
      & while_stage_0_4;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse = PECoreRun_wen & and_dcpl_421
      & (~ accum_vector_operator_1_for_asn_73_itm_2) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2
      & and_dcpl_419;
  assign and_747_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 & reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse;
  assign and_749_cse = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign input_mem_banks_read_read_data_and_33_enex5 = PECoreRun_wen & and_dcpl_421
      & accum_vector_operator_1_for_asn_73_itm_2 & and_dcpl_76 & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo;
  assign mux_95_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, (~ or_tmp_108),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign PECore_DecodeAxiRead_switch_lp_and_23_cse = PECoreRun_wen & mux_95_nl &
      while_stage_0_5;
  assign rva_out_reg_data_and_101_cse = PECoreRun_wen & and_dcpl_434 & (~ accum_vector_operator_1_for_asn_43_itm_2)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 & (~ rva_in_reg_rw_sva_3) &
      (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 | accum_vector_operator_1_for_asn_28_itm_2))
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5 & (~ pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1);
  assign rva_out_reg_data_and_168_enex5 = rva_out_reg_data_and_101_cse & reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_169_enex5 = rva_out_reg_data_and_101_cse & reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_170_enex5 = rva_out_reg_data_and_101_cse & reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_104_cse = PECoreRun_wen & and_dcpl_434 & and_dcpl_419;
  assign rva_out_reg_data_and_171_enex5 = rva_out_reg_data_and_104_cse & reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_172_enex5 = rva_out_reg_data_and_104_cse & reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_173_enex5 = rva_out_reg_data_and_104_cse & reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_174_enex5 = rva_out_reg_data_and_104_cse & reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_175_enex5 = rva_out_reg_data_and_104_cse & reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse = PECoreRun_wen & and_dcpl_445
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 & and_dcpl_155;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse = PECoreRun_wen & and_dcpl_445
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign input_mem_banks_read_read_data_and_34_enex5 = PECoreRun_wen & and_dcpl_415
      & accum_vector_operator_1_for_asn_73_itm_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1;
  assign rva_out_reg_data_and_109_cse = PECoreRun_wen & (~(accum_vector_operator_1_for_asn_73_itm_1
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_2)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1
      & (~(reg_rva_in_reg_rw_sva_2_cse | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign rva_out_reg_data_and_176_enex5 = rva_out_reg_data_and_109_cse & reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  assign rva_out_reg_data_and_177_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_178_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_179_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_180_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse
      & reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_181_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse
      & reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse = PECoreRun_wen & mux_tmp_95
      & and_dcpl_464;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse = PECoreRun_wen & and_dcpl_464;
  assign PECore_DecodeAxiRead_switch_lp_and_29_cse = PECoreRun_wen & (nor_374_cse
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign rva_out_reg_data_and_117_enex5 = PECoreRun_wen & and_dcpl_477 & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[3:1]==3'b010)
      & (~(reg_rva_in_reg_rw_sva_st_1_1_cse | PECore_DecodeAxiRead_switch_lp_nor_tmp_1
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2)) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_182_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_183_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_184_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_185_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse
      & reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_186_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse
      & reg_pe_config_input_counter_sva_dfm_1_enexo;
  assign PECore_DecodeAxiRead_switch_lp_nor_2_cse = ~((while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[3])
      | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[1])
      | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[0]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse = PECoreRun_wen & (~((~(mux_tmp_95
      & nor_374_cse)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_35_cse = PECoreRun_wen & mux_tmp_95
      & nor_374_cse & (~ PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse = PECoreRun_wen & and_dcpl_218
      & and_dcpl_220 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_40_cse = PECoreRun_wen & and_dcpl_314
      & (~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])))
      & nand_34_cse;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse = PECoreRun_wen & (or_dcpl_146
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]!=2'b10)) & and_dcpl_263;
  assign accum_vector_data_mux_57_nl = MUX_v_31_2_2(accum_vector_data_4_sva_4_mx0w0,
      accum_vector_data_4_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_55_nl = MUX_v_31_2_2(accum_vector_data_4_sva_5_mx0w0,
      accum_vector_data_4_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_53_nl = MUX_v_31_2_2(accum_vector_data_4_sva_6_mx0w0,
      accum_vector_data_4_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_21_nl = accum_vector_data_mux_57_nl + accum_vector_data_mux_55_nl
      + accum_vector_data_mux_53_nl;
  assign accum_vector_data_acc_21_nl = nl_accum_vector_data_acc_21_nl[30:0];
  assign accum_vector_data_mux_51_nl = MUX_v_31_2_2(accum_vector_data_4_sva_7_mx0w0,
      accum_vector_data_4_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_49_nl = MUX_v_31_2_2(accum_vector_data_4_sva_8_mx0w0,
      accum_vector_data_4_sva_8, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_47_nl = MUX_v_31_2_2(accum_vector_data_4_sva_9_mx0w0,
      accum_vector_data_4_sva_9, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_22_nl = accum_vector_data_mux_51_nl + accum_vector_data_mux_49_nl
      + accum_vector_data_mux_47_nl;
  assign accum_vector_data_acc_22_nl = nl_accum_vector_data_acc_22_nl[30:0];
  assign nl_accum_vector_data_acc_20_itm = accum_vector_data_acc_21_nl + accum_vector_data_acc_22_nl;
  assign accum_vector_data_acc_20_itm = nl_accum_vector_data_acc_20_itm[30:0];
  assign accum_vector_data_mux_79_nl = MUX_v_31_2_2(accum_vector_data_2_sva_4_mx0w0,
      accum_vector_data_2_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_77_nl = MUX_v_31_2_2(accum_vector_data_2_sva_5_mx0w0,
      accum_vector_data_2_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_75_nl = MUX_v_31_2_2(accum_vector_data_2_sva_6_mx0w0,
      accum_vector_data_2_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_15_nl = accum_vector_data_mux_79_nl + accum_vector_data_mux_77_nl
      + accum_vector_data_mux_75_nl;
  assign accum_vector_data_acc_15_nl = nl_accum_vector_data_acc_15_nl[30:0];
  assign accum_vector_data_mux_73_nl = MUX_v_31_2_2(accum_vector_data_2_sva_7_mx0w0,
      accum_vector_data_2_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_71_nl = MUX_v_31_2_2(accum_vector_data_2_sva_8_mx0w0,
      accum_vector_data_2_sva_8, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_69_nl = MUX_v_31_2_2(accum_vector_data_2_sva_9_mx0w0,
      accum_vector_data_2_sva_9, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_16_nl = accum_vector_data_mux_73_nl + accum_vector_data_mux_71_nl
      + accum_vector_data_mux_69_nl;
  assign accum_vector_data_acc_16_nl = nl_accum_vector_data_acc_16_nl[30:0];
  assign nl_accum_vector_data_acc_14_itm = accum_vector_data_acc_15_nl + accum_vector_data_acc_16_nl;
  assign accum_vector_data_acc_14_itm = nl_accum_vector_data_acc_14_itm[30:0];
  assign accum_vector_data_mux_45_nl = MUX_v_31_2_2(accum_vector_data_5_sva_4_mx0w0,
      accum_vector_data_5_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_43_nl = MUX_v_31_2_2(accum_vector_data_5_sva_5_mx0w0,
      accum_vector_data_5_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_41_nl = MUX_v_31_2_2(accum_vector_data_5_sva_6_mx0w0,
      accum_vector_data_5_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_24_nl = accum_vector_data_mux_45_nl + accum_vector_data_mux_43_nl
      + accum_vector_data_mux_41_nl;
  assign accum_vector_data_acc_24_nl = nl_accum_vector_data_acc_24_nl[30:0];
  assign accum_vector_data_mux_39_nl = MUX_v_31_2_2(accum_vector_data_5_sva_7_mx0w0,
      accum_vector_data_5_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_37_nl = MUX_v_31_2_2(accum_vector_data_5_sva_8_mx0w0,
      accum_vector_data_5_sva_8, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_25_nl = accum_vector_data_mux_39_nl + accum_vector_data_mux_37_nl
      + accum_vector_data_5_sva_9;
  assign accum_vector_data_acc_25_nl = nl_accum_vector_data_acc_25_nl[30:0];
  assign nl_accum_vector_data_acc_23_itm = accum_vector_data_acc_24_nl + accum_vector_data_acc_25_nl;
  assign accum_vector_data_acc_23_itm = nl_accum_vector_data_acc_23_itm[30:0];
  assign accum_vector_data_mux_89_nl = MUX_v_31_2_2(accum_vector_data_1_sva_4_mx0w0,
      accum_vector_data_1_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_87_nl = MUX_v_31_2_2(accum_vector_data_1_sva_5_mx0w0,
      accum_vector_data_1_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_85_nl = MUX_v_31_2_2(accum_vector_data_1_sva_6_mx0w0,
      accum_vector_data_1_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_12_nl = accum_vector_data_mux_89_nl + accum_vector_data_mux_87_nl
      + accum_vector_data_mux_85_nl;
  assign accum_vector_data_acc_12_nl = nl_accum_vector_data_acc_12_nl[30:0];
  assign accum_vector_data_mux_83_nl = MUX_v_31_2_2(accum_vector_data_1_sva_7_mx0w0,
      accum_vector_data_1_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_81_nl = MUX_v_31_2_2(accum_vector_data_1_sva_8_mx0w0,
      accum_vector_data_1_sva_8, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_13_nl = accum_vector_data_mux_83_nl + accum_vector_data_mux_81_nl
      + accum_vector_data_1_sva_9;
  assign accum_vector_data_acc_13_nl = nl_accum_vector_data_acc_13_nl[30:0];
  assign nl_accum_vector_data_acc_11_itm = accum_vector_data_acc_12_nl + accum_vector_data_acc_13_nl;
  assign accum_vector_data_acc_11_itm = nl_accum_vector_data_acc_11_itm[30:0];
  assign accum_vector_data_mux_35_nl = MUX_v_31_2_2(accum_vector_data_6_sva_4_mx0w0,
      accum_vector_data_6_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_33_nl = MUX_v_31_2_2(accum_vector_data_6_sva_5_mx0w0,
      accum_vector_data_6_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_31_nl = MUX_v_31_2_2(accum_vector_data_6_sva_6_mx0w0,
      accum_vector_data_6_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_27_nl = accum_vector_data_mux_35_nl + accum_vector_data_mux_33_nl
      + accum_vector_data_mux_31_nl;
  assign accum_vector_data_acc_27_nl = nl_accum_vector_data_acc_27_nl[30:0];
  assign accum_vector_data_mux_29_nl = MUX_v_31_2_2(accum_vector_data_6_sva_7_mx0w0,
      accum_vector_data_6_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_27_nl = MUX_v_31_2_2(accum_vector_data_6_sva_8_mx0w0,
      accum_vector_data_6_sva_8, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_28_nl = accum_vector_data_mux_29_nl + accum_vector_data_mux_27_nl
      + accum_vector_data_6_sva_9;
  assign accum_vector_data_acc_28_nl = nl_accum_vector_data_acc_28_nl[30:0];
  assign nl_accum_vector_data_acc_26_itm = accum_vector_data_acc_27_nl + accum_vector_data_acc_28_nl;
  assign accum_vector_data_acc_26_itm = nl_accum_vector_data_acc_26_itm[30:0];
  assign accum_vector_data_mux_99_nl = MUX_v_31_2_2(accum_vector_data_0_sva_4_mx0w0,
      accum_vector_data_0_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_97_nl = MUX_v_31_2_2(accum_vector_data_0_sva_5_mx0w0,
      accum_vector_data_0_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_95_nl = MUX_v_31_2_2(accum_vector_data_0_sva_6_mx0w0,
      accum_vector_data_0_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_9_nl = accum_vector_data_mux_99_nl + accum_vector_data_mux_97_nl
      + accum_vector_data_mux_95_nl;
  assign accum_vector_data_acc_9_nl = nl_accum_vector_data_acc_9_nl[30:0];
  assign accum_vector_data_mux_93_nl = MUX_v_31_2_2(accum_vector_data_0_sva_7_mx0w0,
      accum_vector_data_0_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_91_nl = MUX_v_31_2_2(accum_vector_data_0_sva_8_mx0w0,
      accum_vector_data_0_sva_8, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_10_nl = accum_vector_data_mux_93_nl + accum_vector_data_mux_91_nl
      + accum_vector_data_0_sva_9;
  assign accum_vector_data_acc_10_nl = nl_accum_vector_data_acc_10_nl[30:0];
  assign nl_accum_vector_data_acc_8_itm = accum_vector_data_acc_9_nl + accum_vector_data_acc_10_nl;
  assign accum_vector_data_acc_8_itm = nl_accum_vector_data_acc_8_itm[30:0];
  assign accum_vector_data_mux_25_nl = MUX_v_31_2_2(accum_vector_data_7_sva_4_mx0w0,
      accum_vector_data_7_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_23_nl = MUX_v_31_2_2(accum_vector_data_7_sva_5_mx0w0,
      accum_vector_data_7_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_21_nl = MUX_v_31_2_2(accum_vector_data_7_sva_6_mx0w0,
      accum_vector_data_7_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_29_nl = accum_vector_data_mux_25_nl + accum_vector_data_mux_23_nl
      + accum_vector_data_mux_21_nl;
  assign accum_vector_data_acc_29_nl = nl_accum_vector_data_acc_29_nl[30:0];
  assign accum_vector_data_mux_19_nl = MUX_v_31_2_2(accum_vector_data_7_sva_7_mx0w0,
      accum_vector_data_7_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_17_nl = MUX_v_31_2_2(accum_vector_data_7_sva_8_mx0w0,
      accum_vector_data_7_sva_8, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_30_nl = accum_vector_data_mux_19_nl + accum_vector_data_mux_17_nl
      + accum_vector_data_7_sva_9;
  assign accum_vector_data_acc_30_nl = nl_accum_vector_data_acc_30_nl[30:0];
  assign nl_accum_vector_data_acc_itm = accum_vector_data_acc_29_nl + accum_vector_data_acc_30_nl;
  assign accum_vector_data_acc_itm = nl_accum_vector_data_acc_itm[30:0];
  assign accum_vector_data_mux_67_nl = MUX_v_31_2_2(accum_vector_data_3_sva_4_mx0w0,
      accum_vector_data_3_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_65_nl = MUX_v_31_2_2(accum_vector_data_3_sva_5_mx0w0,
      accum_vector_data_3_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_63_nl = MUX_v_31_2_2(accum_vector_data_3_sva_6_mx0w0,
      accum_vector_data_3_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_18_nl = accum_vector_data_mux_67_nl + accum_vector_data_mux_65_nl
      + accum_vector_data_mux_63_nl;
  assign accum_vector_data_acc_18_nl = nl_accum_vector_data_acc_18_nl[30:0];
  assign accum_vector_data_mux_61_nl = MUX_v_31_2_2(accum_vector_data_3_sva_7_mx0w0,
      accum_vector_data_3_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_59_nl = MUX_v_31_2_2(accum_vector_data_3_sva_8_mx0w0,
      accum_vector_data_3_sva_8, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_19_nl = accum_vector_data_mux_61_nl + accum_vector_data_mux_59_nl
      + accum_vector_data_3_sva_9;
  assign accum_vector_data_acc_19_nl = nl_accum_vector_data_acc_19_nl[30:0];
  assign nl_accum_vector_data_acc_17_itm = accum_vector_data_acc_18_nl + accum_vector_data_acc_19_nl;
  assign accum_vector_data_acc_17_itm = nl_accum_vector_data_acc_17_itm[30:0];
  assign and_545_cse = while_stage_0_11 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
      & (~ rva_in_reg_rw_sva_st_1_9);
  assign or_407_cse = (state_2_1_sva!=2'b00) | state_0_sva;
  assign and_549_cse = while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)
      & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  assign weight_port_read_out_data_7_1_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]), weight_port_read_out_data_7_1_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_28_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign ProductSum_for_mux_nl = MUX_v_31_2_2(accum_vector_data_7_sva_8, ProductSum_for_acc_19_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_56_nl = ~ accum_vector_operator_1_for_asn_115_itm_7;
  assign accum_vector_data_7_sva_8_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_nl, accum_vector_operator_1_for_not_56_nl);
  assign ProductSum_for_mux_1_nl = MUX_v_31_2_2(accum_vector_data_7_sva_7, ProductSum_for_acc_18_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_57_nl = ~ accum_vector_operator_1_for_asn_115_itm_7;
  assign accum_vector_data_7_sva_7_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_1_nl, accum_vector_operator_1_for_not_57_nl);
  assign ProductSum_for_mux_2_nl = MUX_v_31_2_2(accum_vector_data_7_sva_6, ProductSum_for_acc_17_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_58_nl = ~ accum_vector_operator_1_for_asn_115_itm_7;
  assign accum_vector_data_7_sva_6_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_2_nl, accum_vector_operator_1_for_not_58_nl);
  assign ProductSum_for_mux_3_nl = MUX_v_31_2_2(accum_vector_data_7_sva_5, ProductSum_for_acc_16_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_59_nl = ~ accum_vector_operator_1_for_asn_115_itm_7;
  assign accum_vector_data_7_sva_5_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_3_nl, accum_vector_operator_1_for_not_59_nl);
  assign ProductSum_for_mux_4_nl = MUX_v_31_2_2(accum_vector_data_7_sva_4, ProductSum_for_acc_15_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_40_nl = ~ accum_vector_operator_1_for_asn_115_itm_7;
  assign accum_vector_data_7_sva_4_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_4_nl, accum_vector_operator_1_for_not_40_nl);
  assign ProductSum_for_mux_5_nl = MUX_v_31_2_2(accum_vector_data_6_sva_8, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_60_nl = ~ accum_vector_operator_1_for_asn_100_itm_7;
  assign accum_vector_data_6_sva_8_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_5_nl, accum_vector_operator_1_for_not_60_nl);
  assign ProductSum_for_mux_6_nl = MUX_v_31_2_2(accum_vector_data_6_sva_7, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_61_nl = ~ accum_vector_operator_1_for_asn_100_itm_7;
  assign accum_vector_data_6_sva_7_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_6_nl, accum_vector_operator_1_for_not_61_nl);
  assign ProductSum_for_mux_7_nl = MUX_v_31_2_2(accum_vector_data_6_sva_6, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_62_nl = ~ accum_vector_operator_1_for_asn_100_itm_7;
  assign accum_vector_data_6_sva_6_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_7_nl, accum_vector_operator_1_for_not_62_nl);
  assign ProductSum_for_mux_8_nl = MUX_v_31_2_2(accum_vector_data_6_sva_5, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_63_nl = ~ accum_vector_operator_1_for_asn_100_itm_7;
  assign accum_vector_data_6_sva_5_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_8_nl, accum_vector_operator_1_for_not_63_nl);
  assign ProductSum_for_mux_9_nl = MUX_v_31_2_2(accum_vector_data_6_sva_4, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_42_nl = ~ accum_vector_operator_1_for_asn_100_itm_7;
  assign accum_vector_data_6_sva_4_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_9_nl, accum_vector_operator_1_for_not_42_nl);
  assign ProductSum_for_mux_10_nl = MUX_v_31_2_2(accum_vector_data_5_sva_8, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_64_nl = ~ accum_vector_operator_1_for_asn_85_itm_7;
  assign accum_vector_data_5_sva_8_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_10_nl, accum_vector_operator_1_for_not_64_nl);
  assign ProductSum_for_mux_11_nl = MUX_v_31_2_2(accum_vector_data_5_sva_7, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_65_nl = ~ accum_vector_operator_1_for_asn_85_itm_7;
  assign accum_vector_data_5_sva_7_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_11_nl, accum_vector_operator_1_for_not_65_nl);
  assign ProductSum_for_mux_12_nl = MUX_v_31_2_2(accum_vector_data_5_sva_6, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_66_nl = ~ accum_vector_operator_1_for_asn_85_itm_7;
  assign accum_vector_data_5_sva_6_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_12_nl, accum_vector_operator_1_for_not_66_nl);
  assign ProductSum_for_mux_13_nl = MUX_v_31_2_2(accum_vector_data_5_sva_5, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_67_nl = ~ accum_vector_operator_1_for_asn_85_itm_7;
  assign accum_vector_data_5_sva_5_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_13_nl, accum_vector_operator_1_for_not_67_nl);
  assign ProductSum_for_mux_14_nl = MUX_v_31_2_2(accum_vector_data_5_sva_4, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_44_nl = ~ accum_vector_operator_1_for_asn_85_itm_7;
  assign accum_vector_data_5_sva_4_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_14_nl, accum_vector_operator_1_for_not_44_nl);
  assign ProductSum_for_mux_15_nl = MUX_v_31_2_2(accum_vector_data_4_sva_9, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_68_nl = ~ accum_vector_operator_1_for_asn_73_itm_7;
  assign accum_vector_data_4_sva_9_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_15_nl, accum_vector_operator_1_for_not_68_nl);
  assign ProductSum_for_mux_16_nl = MUX_v_31_2_2(accum_vector_data_4_sva_8, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_69_nl = ~ accum_vector_operator_1_for_asn_73_itm_7;
  assign accum_vector_data_4_sva_8_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_16_nl, accum_vector_operator_1_for_not_69_nl);
  assign ProductSum_for_mux_17_nl = MUX_v_31_2_2(accum_vector_data_4_sva_7, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_70_nl = ~ accum_vector_operator_1_for_asn_73_itm_7;
  assign accum_vector_data_4_sva_7_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_17_nl, accum_vector_operator_1_for_not_70_nl);
  assign ProductSum_for_mux_18_nl = MUX_v_31_2_2(accum_vector_data_4_sva_6, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_71_nl = ~ accum_vector_operator_1_for_asn_73_itm_7;
  assign accum_vector_data_4_sva_6_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_18_nl, accum_vector_operator_1_for_not_71_nl);
  assign ProductSum_for_mux_19_nl = MUX_v_31_2_2(accum_vector_data_4_sva_5, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_72_nl = ~ accum_vector_operator_1_for_asn_73_itm_7;
  assign accum_vector_data_4_sva_5_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_19_nl, accum_vector_operator_1_for_not_72_nl);
  assign ProductSum_for_mux_20_nl = MUX_v_31_2_2(accum_vector_data_4_sva_4, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_46_nl = ~ accum_vector_operator_1_for_asn_73_itm_7;
  assign accum_vector_data_4_sva_4_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_20_nl, accum_vector_operator_1_for_not_46_nl);
  assign ProductSum_for_mux_21_nl = MUX_v_31_2_2(accum_vector_data_3_sva_8, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_73_nl = ~ accum_vector_operator_1_for_asn_55_itm_7;
  assign accum_vector_data_3_sva_8_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_21_nl, accum_vector_operator_1_for_not_73_nl);
  assign ProductSum_for_mux_22_nl = MUX_v_31_2_2(accum_vector_data_3_sva_7, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_74_nl = ~ accum_vector_operator_1_for_asn_55_itm_7;
  assign accum_vector_data_3_sva_7_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_22_nl, accum_vector_operator_1_for_not_74_nl);
  assign ProductSum_for_mux_23_nl = MUX_v_31_2_2(accum_vector_data_3_sva_6, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_75_nl = ~ accum_vector_operator_1_for_asn_55_itm_7;
  assign accum_vector_data_3_sva_6_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_23_nl, accum_vector_operator_1_for_not_75_nl);
  assign ProductSum_for_mux_24_nl = MUX_v_31_2_2(accum_vector_data_3_sva_5, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_76_nl = ~ accum_vector_operator_1_for_asn_55_itm_7;
  assign accum_vector_data_3_sva_5_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_24_nl, accum_vector_operator_1_for_not_76_nl);
  assign ProductSum_for_mux_25_nl = MUX_v_31_2_2(accum_vector_data_3_sva_4, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_48_nl = ~ accum_vector_operator_1_for_asn_55_itm_7;
  assign accum_vector_data_3_sva_4_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_25_nl, accum_vector_operator_1_for_not_48_nl);
  assign ProductSum_for_mux_26_nl = MUX_v_31_2_2(accum_vector_data_2_sva_9, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_77_nl = ~ accum_vector_operator_1_for_asn_43_itm_7;
  assign accum_vector_data_2_sva_9_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_26_nl, accum_vector_operator_1_for_not_77_nl);
  assign ProductSum_for_mux_27_nl = MUX_v_31_2_2(accum_vector_data_2_sva_8, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_78_nl = ~ accum_vector_operator_1_for_asn_43_itm_7;
  assign accum_vector_data_2_sva_8_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_27_nl, accum_vector_operator_1_for_not_78_nl);
  assign ProductSum_for_mux_28_nl = MUX_v_31_2_2(accum_vector_data_2_sva_7, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_79_nl = ~ accum_vector_operator_1_for_asn_43_itm_7;
  assign accum_vector_data_2_sva_7_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_28_nl, accum_vector_operator_1_for_not_79_nl);
  assign ProductSum_for_mux_29_nl = MUX_v_31_2_2(accum_vector_data_2_sva_6, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_80_nl = ~ accum_vector_operator_1_for_asn_43_itm_7;
  assign accum_vector_data_2_sva_6_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_29_nl, accum_vector_operator_1_for_not_80_nl);
  assign ProductSum_for_mux_30_nl = MUX_v_31_2_2(accum_vector_data_2_sva_5, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_81_nl = ~ accum_vector_operator_1_for_asn_43_itm_7;
  assign accum_vector_data_2_sva_5_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_30_nl, accum_vector_operator_1_for_not_81_nl);
  assign ProductSum_for_mux_31_nl = MUX_v_31_2_2(accum_vector_data_2_sva_4, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_50_nl = ~ accum_vector_operator_1_for_asn_43_itm_7;
  assign accum_vector_data_2_sva_4_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_31_nl, accum_vector_operator_1_for_not_50_nl);
  assign ProductSum_for_mux_32_nl = MUX_v_31_2_2(accum_vector_data_1_sva_8, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_82_nl = ~ accum_vector_operator_1_for_asn_25_itm_7;
  assign accum_vector_data_1_sva_8_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_32_nl, accum_vector_operator_1_for_not_82_nl);
  assign ProductSum_for_mux_33_nl = MUX_v_31_2_2(accum_vector_data_1_sva_7, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_83_nl = ~ accum_vector_operator_1_for_asn_25_itm_7;
  assign accum_vector_data_1_sva_7_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_33_nl, accum_vector_operator_1_for_not_83_nl);
  assign ProductSum_for_mux_34_nl = MUX_v_31_2_2(accum_vector_data_1_sva_6, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_84_nl = ~ accum_vector_operator_1_for_asn_25_itm_7;
  assign accum_vector_data_1_sva_6_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_34_nl, accum_vector_operator_1_for_not_84_nl);
  assign ProductSum_for_mux_35_nl = MUX_v_31_2_2(accum_vector_data_1_sva_5, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_85_nl = ~ accum_vector_operator_1_for_asn_25_itm_7;
  assign accum_vector_data_1_sva_5_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_35_nl, accum_vector_operator_1_for_not_85_nl);
  assign ProductSum_for_mux_36_nl = MUX_v_31_2_2(accum_vector_data_1_sva_4, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_52_nl = ~ accum_vector_operator_1_for_asn_25_itm_7;
  assign accum_vector_data_1_sva_4_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_36_nl, accum_vector_operator_1_for_not_52_nl);
  assign ProductSum_for_mux_37_nl = MUX_v_31_2_2(accum_vector_data_0_sva_8, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_86_nl = ~ accum_vector_operator_1_for_asn_10_itm_7;
  assign accum_vector_data_0_sva_8_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_37_nl, accum_vector_operator_1_for_not_86_nl);
  assign ProductSum_for_mux_38_nl = MUX_v_31_2_2(accum_vector_data_0_sva_7, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_87_nl = ~ accum_vector_operator_1_for_asn_10_itm_7;
  assign accum_vector_data_0_sva_7_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_38_nl, accum_vector_operator_1_for_not_87_nl);
  assign ProductSum_for_mux_39_nl = MUX_v_31_2_2(accum_vector_data_0_sva_6, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_88_nl = ~ accum_vector_operator_1_for_asn_10_itm_7;
  assign accum_vector_data_0_sva_6_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_39_nl, accum_vector_operator_1_for_not_88_nl);
  assign ProductSum_for_mux_40_nl = MUX_v_31_2_2(accum_vector_data_0_sva_5, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_89_nl = ~ accum_vector_operator_1_for_asn_10_itm_7;
  assign accum_vector_data_0_sva_5_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_40_nl, accum_vector_operator_1_for_not_89_nl);
  assign ProductSum_for_mux_41_nl = MUX_v_31_2_2(accum_vector_data_0_sva_4, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign accum_vector_operator_1_for_not_54_nl = ~ accum_vector_operator_1_for_asn_10_itm_7;
  assign accum_vector_data_0_sva_4_mx0w0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ProductSum_for_mux_41_nl, accum_vector_operator_1_for_not_54_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_1
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2!=3'b000));
  assign Arbiter_8U_Roundrobin_pick_nand_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1)
      & and_dcpl_82)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_44_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1
      & and_dcpl_82;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_56_nl = weight_mem_read_arbxbar_arbiters_next_7_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_56_nl,
      weight_mem_read_arbxbar_arbiters_next_7_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_57_nl = weight_mem_read_arbxbar_arbiters_next_7_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_57_nl,
      weight_mem_read_arbxbar_arbiters_next_7_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_58_nl = weight_mem_read_arbxbar_arbiters_next_7_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_58_nl,
      weight_mem_read_arbxbar_arbiters_next_7_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_59_nl = weight_mem_read_arbxbar_arbiters_next_7_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_59_nl,
      weight_mem_read_arbxbar_arbiters_next_7_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_60_nl = weight_mem_read_arbxbar_arbiters_next_7_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_60_nl,
      weight_mem_read_arbxbar_arbiters_next_7_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_61_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_61_nl,
      weight_mem_read_arbxbar_arbiters_next_7_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_82);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign Arbiter_8U_Roundrobin_pick_nand_52_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)
      & and_dcpl_82)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_42_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1
      & and_dcpl_82;
  assign weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_52_cse , Arbiter_8U_Roundrobin_pick_and_42_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_52_cse , Arbiter_8U_Roundrobin_pick_and_42_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_52_cse , Arbiter_8U_Roundrobin_pick_and_42_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_52_cse , Arbiter_8U_Roundrobin_pick_and_42_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_52_cse , Arbiter_8U_Roundrobin_pick_and_42_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_52_cse , Arbiter_8U_Roundrobin_pick_and_42_cse});
  assign weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_82);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign Arbiter_8U_Roundrobin_pick_nand_40_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1)
      & and_dcpl_82)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_36_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1
      & and_dcpl_82;
  assign weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_40_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_40_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_39_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_39_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_40_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_38_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_38_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_40_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_37_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_37_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_40_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_40_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_82);
  assign Arbiter_8U_Roundrobin_pick_nand_65_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1)
      & and_dcpl_82)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_56_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1
      & and_dcpl_82;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_74_nl = weight_mem_read_arbxbar_arbiters_next_4_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_74_nl,
      weight_mem_read_arbxbar_arbiters_next_4_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_65_cse , Arbiter_8U_Roundrobin_pick_and_56_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_cse = weight_mem_read_arbxbar_arbiters_next_4_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_cse,
      weight_mem_read_arbxbar_arbiters_next_4_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_65_cse , Arbiter_8U_Roundrobin_pick_and_56_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_65_cse , Arbiter_8U_Roundrobin_pick_and_56_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_65_cse , Arbiter_8U_Roundrobin_pick_and_56_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_65_cse , Arbiter_8U_Roundrobin_pick_and_56_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_65_cse , Arbiter_8U_Roundrobin_pick_and_56_cse});
  assign weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_82);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign Arbiter_8U_Roundrobin_pick_nand_20_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1)
      & and_dcpl_82)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_26_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1
      & and_dcpl_82;
  assign weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_84_nl = weight_mem_read_arbxbar_arbiters_next_3_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_84_nl,
      weight_mem_read_arbxbar_arbiters_next_3_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_85_nl = weight_mem_read_arbxbar_arbiters_next_3_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_85_nl,
      weight_mem_read_arbxbar_arbiters_next_3_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_82);
  assign Arbiter_8U_Roundrobin_pick_nand_74_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1)
      & and_dcpl_82)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_61_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1
      & and_dcpl_82;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl = weight_mem_read_arbxbar_arbiters_next_2_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl,
      weight_mem_read_arbxbar_arbiters_next_2_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_74_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl = weight_mem_read_arbxbar_arbiters_next_2_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl,
      weight_mem_read_arbxbar_arbiters_next_2_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_74_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl = weight_mem_read_arbxbar_arbiters_next_2_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl,
      weight_mem_read_arbxbar_arbiters_next_2_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_74_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl = weight_mem_read_arbxbar_arbiters_next_2_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl,
      weight_mem_read_arbxbar_arbiters_next_2_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_74_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl,
      weight_mem_read_arbxbar_arbiters_next_2_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_74_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl = weight_mem_read_arbxbar_arbiters_next_2_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl,
      weight_mem_read_arbxbar_arbiters_next_2_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_74_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_82);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign Arbiter_8U_Roundrobin_pick_nand_14_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1)
      & and_dcpl_82)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_23_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1
      & and_dcpl_82;
  assign weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_14_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_12_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_12_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_14_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_11_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_11_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_14_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_14_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_9_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign Arbiter_8U_Roundrobin_pick_1_mux_133_mx1w1 = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_9_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_14_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_8_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_8_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_14_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_82);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign Arbiter_8U_Roundrobin_pick_1_mux_63_mx1w1 = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign Arbiter_8U_Roundrobin_pick_or_2_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1)
      & and_dcpl_82)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_5_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1
      & and_dcpl_82;
  assign weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_or_2_cse , Arbiter_8U_Roundrobin_pick_and_5_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign Arbiter_8U_Roundrobin_pick_1_mux_62_mx1w1 = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_or_2_cse , Arbiter_8U_Roundrobin_pick_and_5_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_4_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_4_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_or_2_cse , Arbiter_8U_Roundrobin_pick_and_5_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_3_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_3_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_or_2_cse , Arbiter_8U_Roundrobin_pick_and_5_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl = weight_mem_read_arbxbar_arbiters_next_0_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl,
      weight_mem_read_arbxbar_arbiters_next_0_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_or_2_cse , Arbiter_8U_Roundrobin_pick_and_5_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_or_2_cse , Arbiter_8U_Roundrobin_pick_and_5_cse});
  assign weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_82);
  assign pe_manager_base_weight_sva_mx1_3_0 = MUX_v_4_2_2((pe_manager_base_weight_sva[3:0]),
      (pe_manager_base_weight_sva_dfm_3_1[3:0]), while_stage_0_5);
  assign pe_manager_base_weight_sva_mx2 = MUX_v_15_2_2(pe_manager_base_weight_sva,
      pe_manager_base_weight_sva_dfm_3_1, while_stage_0_5);
  assign pe_manager_base_weight_sva_mx3_0 = MUX_s_1_2_2((pe_manager_base_weight_sva[0]),
      (pe_manager_base_weight_sva_dfm_3_1[0]), while_stage_0_5);
  assign nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000001;
  assign PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_1_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000001;
  assign operator_15_false_acc_nl = nl_operator_15_false_acc_nl[13:0];
  assign weight_read_addrs_2_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000011;
  assign PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_3_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_1_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:2])}) + 13'b0000000000001;
  assign operator_15_false_acc_1_nl = nl_operator_15_false_acc_1_nl[12:0];
  assign weight_read_addrs_4_14_2_lpi_1_dfm_1_1 = MUX_v_13_2_2(13'b0000000000000,
      operator_15_false_acc_1_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000101;
  assign PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_5_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_2_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000011;
  assign operator_15_false_acc_2_nl = nl_operator_15_false_acc_2_nl[13:0];
  assign weight_read_addrs_6_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_2_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000111;
  assign PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_7_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112, and_107_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97, and_114_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82, and_121_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67, and_dcpl_598);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52, and_135_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37, and_142_cse);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_56_tmp & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_56_tmp & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_60_tmp & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22, and_dcpl_619);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7, and_156_cse);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_34_tmp = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_tmp = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  assign accum_vector_data_3_sva_1_load_mx0w1 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_3_sva_1_load;
  assign PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1 = (state_2_1_sva[0]) & (~((state_2_1_sva[1])
      | state_0_sva));
  assign state_mux_1_cse = MUX_v_2_2_2(state_2_1_sva, state_2_1_sva_dfm_1, while_stage_0_3);
  assign state_0_sva_mx1 = MUX_s_1_2_2(PECore_UpdateFSM_next_state_0_lpi_1_dfm_4,
      state_0_sva, or_dcpl_259);
  assign pe_config_manager_counter_sva_mx1 = MUX_v_4_2_2(pe_config_manager_counter_sva,
      pe_config_manager_counter_sva_dfm_3_1, and_1287_cse);
  assign PECore_PushOutput_PECore_PushOutput_if_and_svs_1 = (state_mux_1_cse[1])
      & (~((state_mux_1_cse[0]) | state_0_sva_mx1));
  assign PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1 = ~(PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_407_cse);
  assign pe_config_input_counter_and_cse = while_if_and_tmp_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign while_and_4_cse = PECore_UpdateFSM_switch_lp_equal_tmp_3_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign nl_operator_8_false_acc_nl = pe_config_input_counter_sva + 8'b00000001;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[7:0];
  assign pe_config_UpdateInputCounter_not_nl = ~ pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl = MUX_v_8_2_2(8'b00000000,
      operator_8_false_acc_nl, pe_config_UpdateInputCounter_not_nl);
  assign pe_config_input_counter_nand_nl = ~(while_stage_0_3 & (~(nor_384_cse | while_and_1266_cse_1)));
  assign pe_config_input_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_input_counter_sva,
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl, pe_config_input_counter_sva_dfm_1,
      {pe_config_input_counter_nand_nl , while_and_4_cse , pe_config_input_counter_and_cse});
  assign nl_operator_8_false_1_acc_nl = pe_config_output_counter_sva + 8'b00000001;
  assign operator_8_false_1_acc_nl = nl_operator_8_false_1_acc_nl[7:0];
  assign pe_config_UpdateManagerCounter_if_not_9_nl = ~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl
      = MUX_v_8_2_2(8'b00000000, operator_8_false_1_acc_nl, pe_config_UpdateManagerCounter_if_not_9_nl);
  assign pe_config_output_counter_nand_nl = ~(while_stage_0_3 & (~((~(and_1600_cse
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1266_cse_1)));
  assign while_and_152_nl = and_1600_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign pe_config_output_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_output_counter_sva,
      pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl,
      pe_config_output_counter_sva_dfm_1, {pe_config_output_counter_nand_nl , while_and_152_nl
      , pe_config_input_counter_and_cse});
  assign while_if_and_2_m1c = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & and_dcpl_206;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl
      = pe_config_is_zero_first_sva & (~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1);
  assign while_if_or_nl = (~((~((~ PECore_UpdateFSM_switch_lp_equal_tmp_5_1) & and_dcpl_206))
      & while_stage_0_3)) | ((~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1)
      & while_if_and_2_m1c);
  assign while_if_and_4_nl = pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
      & while_if_and_2_m1c;
  assign pe_config_is_zero_first_sva_mx1 = MUX1HOT_s_1_3_2(while_if_mux_27_itm_1,
      pe_config_is_zero_first_sva, pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl,
      {and_dcpl_205 , while_if_or_nl , while_if_and_4_nl});
  assign PECore_UpdateFSM_switch_lp_equal_tmp_6 = state_0_sva_mx1 & (state_mux_1_cse==2'b00);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1 = (state_mux_1_cse[0])
      & (~((state_mux_1_cse[1]) | state_0_sva_mx1));
  assign pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1
      = ~((pe_config_manager_counter_sva_mx1 != (operator_4_false_acc_sdt_sva_1[3:0]))
      | (operator_4_false_acc_sdt_sva_1[4]));
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0110);
  assign weight_port_read_out_data_0_7_sva_mx0 = MUX1HOT_v_8_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1,
      weight_port_read_out_data_0_7_sva_dfm_1_1, weight_port_read_out_data_0_7_sva,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_5_sva_mx0 = MUX1HOT_v_8_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1,
      weight_port_read_out_data_0_5_sva_dfm_1_1, weight_port_read_out_data_0_5_sva,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp;
  assign weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  assign weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6,
      or_dcpl_258);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0,
      or_dcpl_258);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5,
      or_dcpl_258);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1,
      or_dcpl_258);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4,
      or_dcpl_258);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2,
      or_dcpl_258);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3,
      or_dcpl_258);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_1_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_60_tmp
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0101);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b111)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1 = (pe_manager_base_weight_sva[2:0]==3'b110)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b100)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b010)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b001)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign weight_mem_run_3_for_land_lpi_1_dfm_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_91_tmp | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1);
  assign weight_mem_run_3_for_land_6_lpi_1_dfm_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_75_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_99_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_111_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_123_tmp);
  assign mux1h_11_nl = MUX1HOT_v_8_7_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[63:56]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63:56]),
      weight_port_read_out_data_0_7_sva_mx0, {and_1006_cse , and_1007_cse , and_1008_cse
      , and_1009_cse , and_1010_cse , and_1011_cse , nor_506_cse});
  assign not_2293_nl = ~ or_dcpl;
  assign weight_port_read_out_data_0_7_sva_dfm_mx0w1 = MUX_v_8_2_2(8'b00000000, mux1h_11_nl,
      not_2293_nl);
  assign or_847_tmp = ((pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2) | and_dcpl;
  assign and_1066_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_847_tmp);
  assign and_1067_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_2_cse & (~ or_847_tmp);
  assign and_1068_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      & (~ or_847_tmp);
  assign and_1069_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      & (~ or_847_tmp);
  assign and_1070_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      & (~ or_847_tmp);
  assign and_1071_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      & (~ or_847_tmp);
  assign nor_512_nl = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_847_tmp);
  assign mux1h_12_nl = MUX1HOT_v_8_7_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[47:40]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[47:40]),
      weight_port_read_out_data_0_5_sva_mx0, {and_1066_nl , and_1067_nl , and_1068_nl
      , and_1069_nl , and_1070_nl , and_1071_nl , nor_512_nl});
  assign not_2295_nl = ~ or_847_tmp;
  assign weight_port_read_out_data_0_5_sva_dfm_mx0w1 = MUX_v_8_2_2(8'b00000000, mux1h_12_nl,
      not_2295_nl);
  assign weight_mem_run_3_for_land_1_lpi_1_dfm_1_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2);
  assign nand_41_cse = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
      & rva_in_reg_rw_sva_st_1_6);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1 = MUX_v_3_2_2(3'b000,
      (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0]), weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp = MUX_s_1_8_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1);
  assign PECore_PushAxiRsp_mux_25_nl = MUX_s_1_2_2(reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse,
      PECore_PushAxiRsp_mux_10_itm_1, rva_in_reg_rw_sva_5);
  assign PECore_PushAxiRsp_if_else_mux_10_mx0w2 = MUX_s_1_2_2(PECore_PushAxiRsp_mux_25_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1);
  assign PECore_PushAxiRsp_if_else_mux_23_mx0w2 = MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1);
  assign while_if_while_if_and_27_nl = MUX_v_8_2_2(8'b00000000, rva_out_reg_data_103_96_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_103_96_sva_dfm_4_mx0w0 = MUX1HOT_v_8_3_2(while_if_while_if_and_27_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_28_nl = MUX_v_8_2_2(8'b00000000, rva_out_reg_data_95_88_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_95_88_sva_dfm_4_mx0w0 = MUX1HOT_v_8_3_2(while_if_while_if_and_28_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_30_nl = MUX_v_8_2_2(8'b00000000, rva_out_reg_data_79_72_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_79_72_sva_dfm_4_mx0w0 = MUX1HOT_v_8_3_2(while_if_while_if_and_30_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_31_nl = MUX_v_8_2_2(8'b00000000, rva_out_reg_data_71_64_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_71_64_sva_dfm_4_mx0w0 = MUX1HOT_v_8_3_2(while_if_while_if_and_31_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_63_sva_dfm_6_mx1 = MUX_s_1_2_2(PECore_PushAxiRsp_mux_23_itm_1,
      rva_out_reg_data_63_sva_dfm_6, nand_76_cse);
  assign rva_out_reg_data_55_48_sva_dfm_6_mx1 = MUX_v_8_2_2(rva_out_reg_data_55_48_sva_dfm_4_1,
      rva_out_reg_data_55_48_sva_dfm_6, or_dcpl_309);
  assign rva_out_reg_data_62_56_sva_dfm_6_mx1 = MUX_v_7_2_2(rva_out_reg_data_62_56_sva_dfm_4_1,
      rva_out_reg_data_62_56_sva_dfm_6, or_dcpl_309);
  assign rva_out_reg_data_46_40_sva_dfm_6_mx1 = MUX_v_7_2_2(rva_out_reg_data_46_40_sva_dfm_4_1,
      rva_out_reg_data_46_40_sva_dfm_6, or_dcpl_309);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1 = MUX_v_4_2_2(rva_out_reg_data_39_36_sva_dfm_4_1,
      rva_out_reg_data_39_36_sva_dfm_6, or_dcpl_309);
  assign rva_out_reg_data_35_32_sva_dfm_6_mx1 = MUX_v_4_2_2(rva_out_reg_data_35_32_sva_dfm_4_1,
      rva_out_reg_data_35_32_sva_dfm_6, or_dcpl_309);
  assign while_and_221_rgt = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_225_rgt = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_229_rgt = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_233_rgt = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_237_rgt = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_241_rgt = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_245_rgt = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_249_rgt = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_253_rgt = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_257_rgt = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_261_rgt = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_265_rgt = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_269_rgt = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_273_rgt = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_277_rgt = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_281_rgt = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_285_rgt = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_289_rgt = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_293_rgt = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_297_rgt = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_301_rgt = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_305_rgt = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_309_rgt = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_313_rgt = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_317_rgt = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_321_rgt = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_325_rgt = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_329_rgt = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_333_rgt = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_337_rgt = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_341_rgt = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_345_rgt = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_349_rgt = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_353_rgt = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_357_rgt = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_361_rgt = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_365_rgt = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_369_rgt = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_373_rgt = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_377_rgt = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_381_rgt = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_385_rgt = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_389_rgt = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_393_rgt = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_397_rgt = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_401_rgt = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_405_rgt = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_409_rgt = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_413_rgt = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_417_rgt = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_421_rgt = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_425_rgt = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_429_rgt = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_433_rgt = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_437_rgt = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_441_rgt = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_445_rgt = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_449_rgt = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_453_rgt = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_457_rgt = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_461_rgt = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_465_rgt = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_469_rgt = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_473_rgt = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_477_rgt = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_481_rgt = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_485_rgt = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_489_rgt = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_493_rgt = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_497_rgt = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_501_rgt = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_505_rgt = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_509_rgt = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_513_rgt = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_517_rgt = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_521_rgt = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_525_rgt = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_529_rgt = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_533_rgt = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_537_rgt = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_541_rgt = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_545_rgt = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_549_rgt = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_553_rgt = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_557_rgt = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_561_rgt = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_565_rgt = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_569_rgt = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_573_rgt = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_577_rgt = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_581_rgt = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_585_rgt = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_589_rgt = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_593_rgt = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_597_rgt = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_601_rgt = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_605_rgt = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_609_rgt = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_613_rgt = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_617_rgt = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_621_rgt = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_625_rgt = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_629_rgt = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_633_rgt = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_637_rgt = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_641_rgt = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_645_rgt = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_649_rgt = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_653_rgt = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_657_rgt = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_661_rgt = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_665_rgt = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_669_rgt = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_673_rgt = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_677_rgt = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_681_rgt = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_685_rgt = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_689_rgt = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_693_rgt = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_697_rgt = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_701_rgt = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_705_rgt = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_709_rgt = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_713_rgt = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_717_rgt = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_721_rgt = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_725_rgt = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_729_rgt = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_733_rgt = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_737_rgt = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_741_rgt = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_745_rgt = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_749_rgt = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_753_rgt = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_757_rgt = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_761_rgt = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_765_rgt = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_769_rgt = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_773_rgt = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_777_rgt = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_781_rgt = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_785_rgt = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_789_rgt = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_793_rgt = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_797_rgt = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_801_rgt = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_805_rgt = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_809_rgt = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_813_rgt = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_817_rgt = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_821_rgt = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_825_rgt = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_829_rgt = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_833_rgt = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_837_rgt = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_841_rgt = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_845_rgt = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_849_rgt = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_853_rgt = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_857_rgt = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_861_rgt = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_865_rgt = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_869_rgt = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_873_rgt = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_877_rgt = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_881_rgt = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_885_rgt = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_889_rgt = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_893_rgt = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_897_rgt = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_901_rgt = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_905_rgt = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_909_rgt = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_913_rgt = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_917_rgt = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_921_rgt = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_925_rgt = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_929_rgt = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_933_rgt = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_937_rgt = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_941_rgt = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_945_rgt = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_949_rgt = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_953_rgt = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_957_rgt = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_961_rgt = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_965_rgt = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_969_rgt = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_973_rgt = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_977_rgt = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_981_rgt = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_985_rgt = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_989_rgt = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_993_rgt = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_997_rgt = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1001_rgt = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1005_rgt = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1009_rgt = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1013_rgt = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1017_rgt = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1021_rgt = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1025_rgt = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1029_rgt = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1033_rgt = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1037_rgt = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1041_rgt = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1045_rgt = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1049_rgt = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1053_rgt = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1057_rgt = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1061_rgt = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1065_rgt = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1069_rgt = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1073_rgt = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1077_rgt = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1081_rgt = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1085_rgt = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1089_rgt = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1093_rgt = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1097_rgt = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1101_rgt = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1105_rgt = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1109_rgt = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1113_rgt = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1117_rgt = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1121_rgt = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1125_rgt = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1129_rgt = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1133_rgt = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1137_rgt = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1141_rgt = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1145_rgt = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1149_rgt = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1153_rgt = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1157_rgt = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1161_rgt = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1165_rgt = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1169_rgt = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1173_rgt = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1177_rgt = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1181_rgt = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1185_rgt = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1189_rgt = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1193_rgt = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1197_rgt = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1201_rgt = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1205_rgt = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1209_rgt = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1213_rgt = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1217_rgt = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1221_rgt = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1225_rgt = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1229_rgt = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1233_rgt = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1237_rgt = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1241_rgt = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign accum_vector_data_5_sva_1_load_mx0w0 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_5_sva_1_load;
  assign input_read_req_valid_lpi_1_dfm_1_mx0w2 = PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
      & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign pe_manager_base_input_sva_mx1_7_0 = MUX_v_8_2_2((pe_manager_base_input_sva[7:0]),
      (pe_manager_base_input_sva_dfm_3_1[7:0]), while_stage_0_3);
  assign pe_manager_base_input_sva_mx2 = MUX_v_15_2_2(pe_manager_base_input_sva,
      pe_manager_base_input_sva_dfm_3_1, while_stage_0_3);
  assign accum_vector_data_7_sva_1_load_mx0w1 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_7_sva_1_load;
  assign accum_vector_data_6_sva_1_load_mx0w1 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_6_sva_1_load;
  assign accum_vector_data_1_sva_1_load_mx0w1 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_1_sva_1_load;
  assign accum_vector_data_0_sva_1_load_mx0w1 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_0_sva_1_load;
  assign accum_vector_data_4_sva_1_load_mx0w0 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_4_sva_1_load;
  assign accum_vector_data_2_sva_1_load_mx0w0 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_2_sva_1_load;
  assign PECore_RunScale_PECore_RunScale_if_and_1_svs_1 = (state_mux_1_cse[0]) &
      state_0_sva_mx1 & (~ (state_mux_1_cse[1]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
      & PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_mx0w0
      | and_315_cse);
  assign PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_DecodeAxiRead_switch_lp_nor_9_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 | PECore_DecodeAxiRead_switch_lp_nor_tmp_9);
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1 = ~(input_read_req_valid_lpi_1_dfm_1_9
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0 = MUX_v_128_2_2(weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0 = MUX_v_120_2_2(weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_8,
      (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:8]), weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {weight_mem_run_3_for_5_and_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b100)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_sva_1 | mux_190_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_sva_1 & (~ mux_190_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_sva_1 | mux_209_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_sva_1 & (~ mux_209_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_sva_1) & and_dcpl_672;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_sva_1 & and_dcpl_672;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]),
      {mux_tmp_171 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_sva_1,
      {mux_tmp_171 , (~ mux_190_itm) , (~ mux_209_itm) , and_dcpl_672});
  assign and_968_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  assign or_565_nl = and_968_cse | or_tmp_205;
  assign mux_219_nl = MUX_s_1_2_2(mux_tmp_195, mux_tmp_194, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign mux_220_nl = MUX_s_1_2_2(or_565_nl, mux_219_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl,
      mux_220_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 | mux_232_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 & (~ mux_232_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 | mux_246_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 & (~ mux_246_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1) & and_dcpl_675;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 & and_dcpl_675;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]),
      {mux_tmp_220 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1,
      {mux_tmp_220 , (~ mux_232_itm) , (~ mux_246_itm) , and_dcpl_675});
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  assign mux_255_nl = MUX_s_1_2_2(or_tmp_284, or_tmp_279, while_stage_0_5);
  assign or_612_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | or_tmp_284;
  assign or_607_nl = while_mux_1437_tmp | or_tmp_279;
  assign mux_254_nl = MUX_s_1_2_2(or_612_nl, or_607_nl, while_stage_0_5);
  assign mux_256_nl = MUX_s_1_2_2(mux_255_nl, mux_254_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl,
      mux_256_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 | mux_272_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 & (~ mux_272_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1) & not_tmp_441;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 & not_tmp_441;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1) & and_dcpl_678;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 & and_dcpl_678;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]),
      {mux_tmp_254 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1,
      {mux_tmp_254 , (~ mux_272_itm) , not_tmp_441 , and_dcpl_678});
  assign and_972_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1;
  assign and_976_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]) & while_mux_1430_tmp;
  assign and_975_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) & while_mux_1435_tmp;
  assign and_971_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  assign and_969_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  assign and_970_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  assign and_973_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) & while_mux_1433_tmp;
  assign and_974_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]) & while_mux_1434_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign nor_500_nl = ~(and_969_cse | and_970_cse | and_971_cse | and_972_cse | or_tmp_305);
  assign nor_501_nl = ~(and_973_cse | and_974_cse | and_975_cse | and_976_cse | or_tmp_297);
  assign mux_287_nl = MUX_s_1_2_2(nor_500_nl, nor_501_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl,
      mux_287_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1) & and_dcpl_679;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 & and_dcpl_679;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1) & and_dcpl_680;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 & and_dcpl_680;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1) & and_dcpl_684;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 & and_dcpl_684;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]),
      {or_dcpl_320 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1,
      operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1, {or_dcpl_320 , and_dcpl_679
      , and_dcpl_680 , and_dcpl_684});
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign mux_322_nl = MUX_s_1_2_2(or_tmp_379, or_tmp_377, while_stage_0_5);
  assign or_708_nl = weight_mem_read_arbxbar_arbiters_next_4_5_sva | or_tmp_379;
  assign or_706_nl = while_mux_1425_tmp | or_tmp_377;
  assign mux_321_nl = MUX_s_1_2_2(or_708_nl, or_706_nl, while_stage_0_5);
  assign mux_323_nl = MUX_s_1_2_2(mux_322_nl, mux_321_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign nor_502_nl = ~(mux_323_nl | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl,
      nor_502_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_24_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1) & and_dcpl_688;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 & and_dcpl_688;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1) & and_dcpl_689;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 & and_dcpl_689;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1) & and_dcpl_695;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 & and_dcpl_695;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]),
      {weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_24_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1,
      operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1, {weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse
      , and_dcpl_688 , and_dcpl_689 , and_dcpl_695});
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse
      = weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign and_709_nl = (~ mux_tmp_323) & and_dcpl_687;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse,
      weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl,
      and_709_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 | mux_340_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 & (~ mux_340_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 | mux_351_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 & (~ mux_351_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1) & and_dcpl_697;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 & and_dcpl_697;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]),
      {mux_tmp_333 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1,
      {mux_tmp_333 , (~ mux_340_itm) , (~ mux_351_itm) , and_dcpl_697});
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  assign mux_359_nl = MUX_s_1_2_2(or_tmp_419, mux_tmp_338, while_stage_0_5);
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, mux_tmp_339, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl,
      mux_360_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 | mux_378_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 & (~ mux_378_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1) & not_tmp_470;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 & not_tmp_470;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1) & and_dcpl_700;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 & and_dcpl_700;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]),
      {mux_tmp_364 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1,
      {mux_tmp_364 , (~ mux_378_itm) , not_tmp_470 , and_dcpl_700});
  assign and_979_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1;
  assign and_978_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]) & weight_mem_read_arbxbar_arbiters_next_0_3_sva;
  assign and_977_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) & weight_mem_read_arbxbar_arbiters_next_0_4_sva;
  assign and_981_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]) & while_mux_1399_tmp;
  assign and_980_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) & while_mux_1398_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign nor_503_nl = ~(and_977_cse | and_978_cse | and_979_cse | or_tmp_460);
  assign mux_396_nl = MUX_s_1_2_2(or_tmp_450, or_tmp_447, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_397_nl = MUX_s_1_2_2(mux_396_nl, mux_tmp_376, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign nor_504_nl = ~(and_980_cse | and_981_cse | mux_397_nl);
  assign mux_398_nl = MUX_s_1_2_2(nor_503_nl, nor_504_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl,
      mux_398_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_123_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_111_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_99_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_91_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_75_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = (pe_manager_base_weight_sva_mx2[14:4])
      + PEManager_15U_GetWeightAddr_else_acc_3_1;
  assign PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1[10:0];
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_1_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_1_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1 | (weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1 | (weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1) & and_dcpl_704;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 & and_dcpl_704;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_44_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1) & and_dcpl_705;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 & and_dcpl_705;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_46_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1) & and_dcpl_708;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_47_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 & and_dcpl_708;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]),
      {weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_44_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_46_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_47_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1,
      operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1, {weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse
      , and_dcpl_704 , and_dcpl_705 , and_dcpl_708});
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse
      = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      = MUX_s_1_2_2(or_222_cse, weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse,
      weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp);
  assign operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp
      = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 | (weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1 | (weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1 | (weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1 | (weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 | (weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]));
  assign operator_7_false_1_operator_7_false_1_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 | (weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]));
  assign weight_read_addrs_0_3_0_lpi_1_dfm_4 = MUX_v_4_2_2(4'b0000, pe_manager_base_weight_sva_mx1_3_0,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_4_false_acc_sdt_sva_1 = conv_u2s_4_5(pe_config_num_manager_sva)
      + 5'b11111;
  assign operator_4_false_acc_sdt_sva_1 = nl_operator_4_false_acc_sdt_sva_1[4:0];
  assign while_and_1266_cse_1 = (~ while_if_and_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_if_and_tmp_1 = PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      = ~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl = start_PopNB_mioi_data_rsc_z_mxwt
      & pe_config_is_valid_sva & start_PopNB_mioi_return_rsc_z_mxwt;
  assign PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl = pe_config_is_zero_first_sva
      & pe_manager_zero_active_sva;
  assign PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl = ~(pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign PECore_UpdateFSM_switch_lp_mux1h_14_nl = MUX1HOT_s_1_4_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl,
      PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl, pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1,
      PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl, {PECore_UpdateFSM_switch_lp_and_7_itm_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_2_1 , PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_5_1});
  assign PECore_UpdateFSM_next_state_0_lpi_1_dfm_4 = PECore_UpdateFSM_switch_lp_mux1h_14_nl
      & PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  assign pe_config_UpdateManagerCounter_if_if_unequal_tmp = pe_config_output_counter_sva
      != (operator_8_false_acc_sdt_sva_1[7:0]);
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      = ~(pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]));
  assign input_write_req_valid_lpi_1_dfm_5 = PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      & PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1 = ~(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign weight_mem_banks_load_store_1_for_else_else_and_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_or_nl = (weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1);
  assign weight_mem_banks_load_store_1_for_else_else_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9 = MUX1HOT_v_8_6_2(BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8,
      ({weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7_4
      , weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_3_0}),
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1,
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[7:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[7:0]),
      {weight_mem_banks_load_store_1_for_else_else_and_nl , weight_mem_banks_load_store_1_for_else_else_or_nl
      , weight_mem_banks_load_store_1_for_else_else_and_4_nl , weight_mem_banks_load_store_1_for_else_else_and_6_nl
      , weight_mem_banks_load_store_1_for_else_else_and_8_nl , weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse = reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_weight_mem_run_3_for_5_and_14_itm_1_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_weight_mem_run_3_for_5_and_14_itm_1_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_265_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_265_nl , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1 , PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {weight_mem_run_3_for_5_and_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {weight_mem_run_3_for_5_and_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {weight_mem_run_3_for_5_and_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {weight_mem_run_3_for_5_and_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {weight_mem_run_3_for_5_and_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_21_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_21_nl
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {weight_mem_run_3_for_5_and_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_nl
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {weight_mem_run_3_for_5_and_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1 = (~(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0,
      or_dcpl_328);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4, nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0,
      or_dcpl_328);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5, nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0,
      or_dcpl_328);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6, nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0,
      or_dcpl_328);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0,
      or_dcpl_328);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0,
      or_dcpl_328);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0,
      or_dcpl_328);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_56_tmp = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_60_tmp = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1 = and_315_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0;
  assign nl_operator_16_false_acc_sdt_sva_1 = conv_u2s_8_9(pe_manager_num_input_sva)
      + 9'b111111111;
  assign operator_16_false_acc_sdt_sva_1 = nl_operator_16_false_acc_sdt_sva_1[8:0];
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1 = ~((state_mux_1_cse!=2'b00)
      | state_0_sva_mx1);
  assign PECore_UpdateFSM_switch_lp_nor_tmp_1 = ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_6 | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1
      | PECore_RunScale_PECore_RunScale_if_and_1_svs_1 | PECore_PushOutput_PECore_PushOutput_if_and_svs_1);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_148_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_108_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[103:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_148_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_163_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_124_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[103:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_163_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_sva_1
      = MUX_v_8_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_108_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_124_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_149_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_107_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[95:88]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_149_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_164_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_123_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[95:88]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_164_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1
      = MUX_v_8_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_107_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_123_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_151_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_102_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[55:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_151_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_166_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_118_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[55:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_166_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_sva_1
      = MUX_v_8_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_102_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_118_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_152_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_105_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[79:72]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_152_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_167_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_121_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[79:72]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_167_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_sva_1
      = MUX_v_8_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_105_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_121_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_153_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_104_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[71:64]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_153_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_168_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_120_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[71:64]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_168_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_sva_1
      = MUX_v_8_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_104_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_120_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign while_and_40_tmp = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp
      = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2) | reg_rva_in_reg_rw_sva_2_cse
      | (~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp!=8'b00000000))) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7])));
  assign PECore_DecodeAxiWrite_switch_lp_or_5_cse_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  assign rva_out_reg_data_63_sva_dfm_7 = rva_out_reg_data_63_sva_dfm_6_mx1 & rva_in_reg_rw_sva_5;
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_1_0_sva_1 = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]!=2'b00));
  assign input_mem_banks_write_if_for_if_and_stg_1_1_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b01);
  assign input_mem_banks_write_if_for_if_and_stg_1_2_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b10);
  assign input_mem_banks_write_if_for_if_and_stg_1_3_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b11);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign nl_PEManager_15U_GetInputAddr_acc_nl = input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt
      + (pe_manager_base_input_sva[7:0]);
  assign PEManager_15U_GetInputAddr_acc_nl = nl_PEManager_15U_GetInputAddr_acc_nl[7:0];
  assign input_write_addrs_lpi_1_dfm_2 = PEManager_15U_GetInputAddr_acc_nl & ({{7{PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1}},
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1})
      & ({{7{PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1}}, PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1});
  assign input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1 = ~((input_write_addrs_lpi_1_dfm_2[1:0]!=2'b00));
  assign input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b01);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b10);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b11);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2
      | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_4 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0011);
  assign PECore_DecodeAxiRead_switch_lp_nor_13_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_not_185 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 =
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:1]!=15'b000000000000000));
  assign PECore_PushAxiRsp_if_asn_79 = (~ rva_in_reg_rw_sva_9) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_81 = rva_in_reg_rw_sva_9 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_83 = input_read_req_valid_lpi_1_dfm_1_9 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign weight_mem_run_3_for_5_asn_447 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_449 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_451 = (weight_read_addrs_7_lpi_1_dfm_3_2_0[2])
      & nor_573_cse & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_453 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_414 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_416 = (weight_read_addrs_5_lpi_1_dfm_3_2_0[2])
      & nor_582_cse & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_418 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_434 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign while_while_nor_259_cse = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_3 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign while_and_39_cse = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign while_and_1243_cse = weight_mem_run_3_for_land_1_lpi_1_dfm_3 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign PECore_PushAxiRsp_if_asn_87 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign PECore_PushAxiRsp_if_asn_89 = (~ rva_in_reg_rw_sva_5) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign PECore_PushAxiRsp_if_asn_91 = rva_in_reg_rw_sva_5 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign while_asn_998 = rva_in_reg_rw_sva_5 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_44_itm_1
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_14_itm_1
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_152 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_156 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_2
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_30_itm_2
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_2
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign Arbiter_8U_Roundrobin_pick_1_mux_589_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1443_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_589_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_590_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1442_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_590_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_591_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1441_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_591_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_592_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1440_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_592_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_593_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1439_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_593_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_594_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1438_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_594_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1437_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_595_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1436_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_595_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_596_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1435_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_596_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_597_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1434_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_597_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_39_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_598_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1433_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_598_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_38_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_599_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1432_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_599_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_37_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_600_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1431_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_600_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1430_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_603_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1427_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_603_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_604_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1426_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_604_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_605_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1425_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_605_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_606_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1424_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_606_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_607_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1422_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_607_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_608_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1421_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_608_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_609_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1420_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_609_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_619_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1408_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_619_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_620_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1407_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_620_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_12_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_621_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1406_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_621_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_11_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_622_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1405_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_622_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_624_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1403_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_624_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_8_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1401_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_63_mx1w1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1400_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_62_mx1w1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_627_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1399_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_627_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_4_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_628_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1398_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_628_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_3_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_630_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1396_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_630_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_dcpl_6 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
      & while_stage_0_10;
  assign and_dcpl_7 = and_dcpl_6 & (~ rva_in_reg_rw_sva_st_1_8);
  assign and_dcpl_8 = and_dcpl_7 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6
      | rva_in_reg_rw_sva_8 | input_read_req_valid_lpi_1_dfm_1_8));
  assign and_dcpl_24 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & while_stage_0_10;
  assign and_dcpl_29 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & while_stage_0_9;
  assign or_tmp_8 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  assign and_cse = rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign and_dcpl_33 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      & while_stage_0_8;
  assign and_dcpl_35 = PECore_RunMac_PECore_RunMac_if_and_svs_st_5 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7;
  assign or_tmp_14 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | rva_in_reg_rw_sva_st_1_5;
  assign or_tmp_15 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_5);
  assign and_dcpl_40 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7;
  assign not_tmp_33 = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_5);
  assign nor_tmp_2 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign or_36_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign mux_15_itm = MUX_s_1_2_2(nor_tmp_2, or_36_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_2);
  assign and_dcpl_47 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7;
  assign and_dcpl_54 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign and_dcpl_55 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign or_tmp_23 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      | rva_in_reg_rw_sva_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1
      | rva_in_reg_rw_sva_st_1_4;
  assign and_tmp_1 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & or_tmp_23;
  assign or_tmp_24 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 | rva_in_reg_rw_sva_4
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 | rva_in_reg_rw_sva_st_1_4;
  assign or_dcpl_12 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ while_stage_0_6);
  assign and_dcpl_76 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_dcpl_82 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_84 = (((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1)
      & and_dcpl_82;
  assign and_dcpl_86 = (((Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 |
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1) | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1)
      & and_dcpl_82;
  assign and_dcpl_88 = (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1
      | and_745_cse | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp)
      & and_dcpl_82;
  assign or_dcpl_41 = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1;
  assign or_85_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp
      | (or_dcpl_41 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1) | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  assign and_dcpl_90 = or_85_cse & and_dcpl_82;
  assign or_dcpl_48 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse;
  assign or_92_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1
      | (or_dcpl_48 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1) | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp;
  assign and_dcpl_92 = or_92_cse & and_dcpl_82;
  assign and_dcpl_94 = (((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1) | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp)
      & and_dcpl_82;
  assign or_106_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1
      | ((Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1) | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_91_tmp;
  assign and_dcpl_96 = or_106_cse & and_dcpl_82;
  assign or_113_cse = ((Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 |
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1) | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_99_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp;
  assign and_dcpl_98 = or_113_cse & and_dcpl_82;
  assign nor_285_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]));
  assign and_107_cse = (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) |
      (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]))) & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]))) & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]))) & nor_285_cse;
  assign nor_286_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]));
  assign and_114_cse = nor_286_cse & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])));
  assign nor_290_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]));
  assign and_121_cse = nor_290_cse & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])));
  assign nor_294_cse = ~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]));
  assign nor_297_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]));
  assign and_135_cse = (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) |
      (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])));
  assign nor_302_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]));
  assign and_142_cse = nor_302_cse & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])));
  assign nor_308_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]));
  assign nor_309_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]));
  assign nor_306_cse = ~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]));
  assign nor_307_cse = ~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]));
  assign nor_310_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]));
  assign and_156_cse = nor_310_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])));
  assign and_dcpl_155 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_162 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign and_dcpl_171 = and_dcpl_155 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]);
  assign and_dcpl_174 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]));
  assign and_dcpl_175 = and_dcpl_155 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]);
  assign and_dcpl_177 = and_dcpl_155 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]))
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign and_dcpl_178 = and_dcpl_155 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]);
  assign and_dcpl_181 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]));
  assign and_dcpl_182 = and_dcpl_155 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]);
  assign and_dcpl_185 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]));
  assign and_dcpl_187 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]) & while_stage_0_4;
  assign and_dcpl_190 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])) & while_stage_0_4;
  assign and_dcpl_191 = and_dcpl_155 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]);
  assign and_dcpl_194 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]));
  assign and_dcpl_196 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_198 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6])
      & and_dcpl_155;
  assign and_dcpl_200 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_202 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7])
      & and_dcpl_155;
  assign and_dcpl_205 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign and_dcpl_206 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign and_dcpl_209 = (state_2_1_sva==2'b01) & (~ state_0_sva) & and_dcpl_206;
  assign mux_26_nl = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      state_2_1_sva[1]);
  assign and_735_nl = (state_2_1_sva[1]) & PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  assign mux_27_nl = MUX_s_1_2_2(mux_26_nl, and_735_nl, state_2_1_sva[0]);
  assign mux_28_nl = MUX_s_1_2_2(mux_27_nl, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      state_0_sva);
  assign and_dcpl_212 = mux_28_nl & (~(PECore_RunFSM_switch_lp_nor_tmp_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign and_dcpl_213 = (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign or_dcpl_146 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]!=2'b01);
  assign and_dcpl_214 = reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign and_dcpl_218 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign and_dcpl_219 = and_dcpl_218 & and_dcpl_214 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_220 = reg_rva_in_PopNB_mioi_iswt0_cse & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_222 = and_dcpl_218 & and_dcpl_220 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_224 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & (~ rva_in_reg_rw_sva_st_1_7);
  assign or_tmp_36 = rva_in_reg_rw_sva_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1
      | rva_in_reg_rw_sva_st_1_4;
  assign or_tmp_37 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      | (~ or_tmp_36);
  assign and_dcpl_248 = PECore_RunFSM_switch_lp_equal_tmp_1_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_736_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  assign or_230_nl = (~ Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1)
      | (~ (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])) | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp;
  assign mux_tmp_42 = MUX_s_1_2_2(or_230_nl, Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp,
      and_736_cse);
  assign mux_tmp_43 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp,
      mux_tmp_42, and_743_cse);
  assign and_738_cse = weight_mem_read_arbxbar_arbiters_next_1_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign or_232_nl = (~(and_738_cse | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]))) | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp;
  assign mux_tmp_47 = MUX_s_1_2_2(or_232_nl, Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp,
      weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign mux_51_nl = MUX_s_1_2_2(mux_tmp_47, mux_tmp_42, weight_mem_read_arbxbar_arbiters_next_1_4_sva);
  assign mux_tmp_49 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp,
      mux_51_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign and_dcpl_262 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
      & while_stage_0_8;
  assign and_dcpl_263 = and_cse & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_277 = and_dcpl_224 & while_stage_0_9;
  assign and_dcpl_284 = (PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 | (~
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7)) & and_dcpl_29;
  assign and_dcpl_290 = and_dcpl_224 & (~ rva_in_reg_rw_sva_7);
  assign and_dcpl_314 = nor_524_cse & and_cse;
  assign and_dcpl_323 = PECore_RunMac_PECore_RunMac_if_and_svs_st_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign and_dcpl_352 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
      & (~ rva_in_reg_rw_sva_st_1_6);
  assign and_dcpl_353 = and_dcpl_352 & while_stage_0_8;
  assign and_dcpl_356 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4
      | rva_in_reg_rw_sva_6 | input_read_req_valid_lpi_1_dfm_1_6);
  assign and_dcpl_382 = while_stage_0_7 & (~ rva_in_reg_rw_sva_st_1_5) & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign or_tmp_85 = PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_5);
  assign or_dcpl_216 = (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp)
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp;
  assign and_dcpl_415 = or_dcpl_216 & (~ reg_rva_in_reg_rw_sva_2_cse);
  assign nor_329_cse = ~(accum_vector_operator_1_for_asn_73_itm_1 | reg_rva_in_reg_rw_sva_2_cse);
  assign and_dcpl_419 = (~ rva_in_reg_rw_sva_3) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_dcpl_421 = ~(pe_manager_base_weight_slc_pe_manager_base_weight_2_0_371_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1);
  assign or_tmp_108 = rva_in_reg_rw_sva_3 | accum_vector_operator_1_for_asn_73_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_371_itm_1;
  assign and_dcpl_434 = and_dcpl_421 & (~ accum_vector_operator_1_for_asn_73_itm_2);
  assign and_dcpl_445 = or_dcpl_216 & nor_329_cse;
  assign or_tmp_112 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 | (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1)));
  assign not_tmp_248 = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 | (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1));
  assign and_dcpl_464 = nor_374_cse & and_dcpl_205;
  assign mux_tmp_95 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1!=4'b0100));
  assign and_dcpl_477 = nor_374_cse & (~(reg_rva_in_reg_rw_sva_st_1_1_cse | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[0])));
  assign and_dcpl_497 = ((~ PECore_UpdateFSM_switch_lp_equal_tmp_2_1) | PECore_UpdateFSM_switch_lp_equal_tmp_5_1)
      & and_dcpl_206;
  assign nand_34_cse = ~(PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]));
  assign and_dcpl_507 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_6 & while_stage_0_8;
  assign and_dcpl_514 = and_dcpl_76 & ProductSum_for_asn_69_itm_3;
  assign or_357_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1;
  assign mux_99_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      or_357_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_tmp_4 = while_stage_0_6 & mux_99_nl;
  assign and_dcpl_516 = and_dcpl_76 & ProductSum_for_asn_56_itm_3;
  assign or_361_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1;
  assign mux_102_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      or_361_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_tmp_5 = while_stage_0_6 & mux_102_nl;
  assign or_365_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
      | ProductSum_for_asn_41_itm_3;
  assign mux_105_nl = MUX_s_1_2_2(or_113_cse, or_365_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_6 = while_stage_0_5 & mux_105_nl;
  assign or_373_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 | ProductSum_for_asn_28_itm_3;
  assign mux_108_nl = MUX_s_1_2_2(or_106_cse, or_373_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_7 = while_stage_0_5 & mux_108_nl;
  assign or_381_nl = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp;
  assign or_380_nl = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp;
  assign mux_tmp_108 = MUX_s_1_2_2(or_381_nl, or_380_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign or_379_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_3 | ProductSum_for_asn_128_itm_3;
  assign mux_112_nl = MUX_s_1_2_2(mux_tmp_108, or_379_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_8 = while_stage_0_5 & mux_112_nl;
  assign or_385_nl = PECore_RunMac_PECore_RunMac_if_and_svs_st_3 | ProductSum_for_asn_108_itm_3;
  assign mux_115_nl = MUX_s_1_2_2(or_92_cse, or_385_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_9 = while_stage_0_5 & mux_115_nl;
  assign or_391_nl = PECore_RunMac_PECore_RunMac_if_and_svs_3 | PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
  assign mux_118_nl = MUX_s_1_2_2(or_85_cse, or_391_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_10 = while_stage_0_5 & mux_118_nl;
  assign or_398_nl = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp;
  assign or_397_nl = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp;
  assign mux_tmp_118 = MUX_s_1_2_2(or_398_nl, or_397_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign or_396_nl = PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 | PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign mux_122_nl = MUX_s_1_2_2(mux_tmp_118, or_396_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_11 = while_stage_0_5 & mux_122_nl;
  assign and_754_cse = PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign and_dcpl_539 = fsm_output & (~ weight_mem_run_3_for_land_3_lpi_1_dfm_3);
  assign and_dcpl_541 = fsm_output & (~ weight_mem_run_3_for_land_5_lpi_1_dfm_3);
  assign and_dcpl_552 = weight_mem_run_3_for_land_7_lpi_1_dfm_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_dcpl_553 = ~(weight_mem_run_3_for_land_7_lpi_1_dfm_2 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_dcpl_243 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
      | (~ while_stage_0_8);
  assign or_dcpl_249 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6);
  assign or_dcpl_251 = (~ weight_mem_run_3_for_land_7_lpi_1_dfm_2) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7);
  assign or_dcpl_252 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7);
  assign or_dcpl_253 = or_dcpl_252 | (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign or_dcpl_255 = or_dcpl_252 | (~ weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign and_dcpl_576 = and_dcpl_82 & (~ while_stage_0_4);
  assign or_dcpl_258 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ while_stage_0_5);
  assign and_dcpl_593 = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) |
      (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]));
  assign and_dcpl_598 = nor_294_cse & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]))) & and_dcpl_593 & nor_297_cse;
  assign and_dcpl_615 = nor_308_cse & nor_309_cse;
  assign and_dcpl_619 = nor_306_cse & nor_307_cse & and_dcpl_615;
  assign or_dcpl_259 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ while_stage_0_3);
  assign or_dcpl_270 = nand_91_cse | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_271 = or_dcpl_146 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]);
  assign and_dcpl_631 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign and_dcpl_632 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]));
  assign and_dcpl_633 = and_dcpl_632 & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign and_dcpl_634 = and_dcpl_632 & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]));
  assign or_dcpl_305 = (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | nand_34_cse;
  assign and_dcpl_637 = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]==2'b10);
  assign and_dcpl_638 = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]!=2'b00));
  assign or_dcpl_309 = nand_76_cse | rva_in_reg_rw_sva_6;
  assign and_dcpl_658 = (~(rva_in_PopNB_mioi_return_rsc_z_mxwt | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign and_dcpl_659 = or_dcpl_259 & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign or_494_nl = while_stage_0_3 | (state_2_1_sva!=2'b01) | state_0_sva;
  assign or_493_nl = (state_2_1_sva!=2'b01) | state_0_sva;
  assign mux_159_nl = MUX_s_1_2_2(or_493_nl, mux_136_cse, while_stage_0_3);
  assign nor_35_nl = ~((state_2_1_sva_dfm_1!=2'b01));
  assign mux_160_nl = MUX_s_1_2_2(or_494_nl, mux_159_nl, nor_35_nl);
  assign and_dcpl_663 = (~ mux_160_nl) & and_dcpl_213;
  assign and_763_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_6_sva;
  assign or_tmp_187 = and_763_cse | (weight_mem_read_arbxbar_arbiters_next_7_5_sva
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]));
  assign or_513_nl = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign mux_tmp_166 = MUX_s_1_2_2(or_tmp_187, or_513_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign and_765_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) & Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1;
  assign or_516_cse = and_765_cse | (Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 &
      (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]));
  assign mux_tmp_167 = MUX_s_1_2_2(or_tmp_187, or_516_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_518_nl = and_968_cse | or_tmp_187;
  assign mux_172_nl = MUX_s_1_2_2(mux_tmp_167, mux_tmp_166, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_517_nl = Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 | mux_tmp_167;
  assign or_515_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | mux_tmp_166;
  assign mux_171_nl = MUX_s_1_2_2(or_517_nl, or_515_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_173_nl = MUX_s_1_2_2(mux_172_nl, mux_171_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign mux_tmp_171 = MUX_s_1_2_2(or_518_nl, mux_173_nl, while_stage_0_5);
  assign nand_tmp_8 = ~(weight_mem_read_arbxbar_arbiters_next_7_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      & (~ or_tmp_187));
  assign and_772_cse = weight_mem_read_arbxbar_arbiters_next_7_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign and_771_cse = weight_mem_read_arbxbar_arbiters_next_7_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign mux_178_nl = MUX_s_1_2_2(nand_tmp_8, or_tmp_187, and_771_cse);
  assign mux_176_nl = MUX_s_1_2_2(nand_tmp_8, or_tmp_187, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign or_522_nl = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign mux_175_nl = MUX_s_1_2_2(nand_tmp_8, or_tmp_187, or_522_nl);
  assign mux_177_nl = MUX_s_1_2_2(mux_176_nl, mux_175_nl, weight_mem_read_arbxbar_arbiters_next_7_3_sva);
  assign mux_179_nl = MUX_s_1_2_2(mux_178_nl, mux_177_nl, weight_mem_read_arbxbar_arbiters_next_7_2_sva);
  assign mux_tmp_177 = MUX_s_1_2_2(mux_179_nl, or_tmp_187, and_772_cse);
  assign or_520_nl = (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])))
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign mux_tmp_178 = MUX_s_1_2_2(mux_tmp_177, or_520_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign and_778_cse = Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign and_777_cse = Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign and_776_cse = Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nand_9_nl = ~(Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      & (~ or_516_cse));
  assign mux_182_nl = MUX_s_1_2_2(nand_9_nl, or_516_cse, and_776_cse);
  assign mux_183_nl = MUX_s_1_2_2(mux_182_nl, or_516_cse, and_777_cse);
  assign mux_184_nl = MUX_s_1_2_2(mux_183_nl, or_516_cse, and_778_cse);
  assign mux_tmp_182 = MUX_s_1_2_2(mux_tmp_177, mux_184_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign mux_188_nl = MUX_s_1_2_2(mux_tmp_182, mux_tmp_178, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_189_nl = MUX_s_1_2_2(mux_tmp_177, mux_188_nl, while_stage_0_5);
  assign or_526_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | mux_tmp_177;
  assign or_525_nl = Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 | mux_tmp_182;
  assign or_523_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | mux_tmp_178;
  assign mux_186_nl = MUX_s_1_2_2(or_525_nl, or_523_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_187_nl = MUX_s_1_2_2(or_526_nl, mux_186_nl, while_stage_0_5);
  assign mux_190_itm = MUX_s_1_2_2(mux_189_nl, mux_187_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign or_tmp_201 = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign nor_tmp_65 = weight_mem_read_arbxbar_arbiters_next_7_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign mux_191_nl = MUX_s_1_2_2((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]),
      or_tmp_201, weight_mem_read_arbxbar_arbiters_next_7_4_sva);
  assign mux_tmp_189 = MUX_s_1_2_2(nor_tmp_65, mux_191_nl, weight_mem_read_arbxbar_arbiters_next_7_5_sva);
  assign and_781_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  assign or_tmp_205 = and_772_cse | and_781_cse | and_771_cse | and_763_cse | mux_tmp_189;
  assign or_527_nl = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign mux_tmp_190 = MUX_s_1_2_2(or_tmp_205, or_527_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign nor_tmp_70 = Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign mux_194_nl = MUX_s_1_2_2((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]),
      or_tmp_201, Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1);
  assign mux_tmp_192 = MUX_s_1_2_2(nor_tmp_70, mux_194_nl, Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1);
  assign or_537_nl = and_778_cse | and_777_cse | and_776_cse | and_765_cse | mux_tmp_192;
  assign mux_tmp_193 = MUX_s_1_2_2(or_tmp_205, or_537_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_538_nl = Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 | mux_tmp_193;
  assign or_533_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | mux_tmp_190;
  assign mux_tmp_194 = MUX_s_1_2_2(or_538_nl, or_533_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_195 = MUX_s_1_2_2(mux_tmp_193, mux_tmp_190, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_213 = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])) |
      (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign mux_199_nl = MUX_s_1_2_2((~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])),
      or_tmp_213, weight_mem_read_arbxbar_arbiters_next_7_4_sva);
  assign or_541_nl = weight_mem_read_arbxbar_arbiters_next_7_5_sva | mux_199_nl;
  assign or_539_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva | mux_tmp_189;
  assign mux_200_nl = MUX_s_1_2_2(or_541_nl, or_539_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign or_tmp_217 = and_772_cse | and_781_cse | and_771_cse | mux_200_nl;
  assign mux_207_nl = MUX_s_1_2_2(or_tmp_217, or_tmp_205, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign or_551_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | or_tmp_205;
  assign mux_208_nl = MUX_s_1_2_2(mux_207_nl, or_551_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign mux_201_nl = MUX_s_1_2_2((~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])),
      or_tmp_213, Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1);
  assign or_547_nl = Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 | mux_201_nl;
  assign or_546_nl = Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 | mux_tmp_192;
  assign mux_202_nl = MUX_s_1_2_2(or_547_nl, or_546_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign or_550_nl = and_778_cse | and_777_cse | and_776_cse | mux_202_nl;
  assign mux_203_nl = MUX_s_1_2_2(or_tmp_217, or_550_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_545_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7])
      | or_tmp_217;
  assign mux_204_nl = MUX_s_1_2_2(mux_203_nl, or_545_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_205_nl = MUX_s_1_2_2(mux_204_nl, mux_tmp_195, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign mux_206_nl = MUX_s_1_2_2(mux_205_nl, mux_tmp_194, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign mux_209_itm = MUX_s_1_2_2(mux_208_nl, mux_206_nl, while_stage_0_5);
  assign or_tmp_225 = and_771_cse | nor_tmp_65;
  assign or_557_nl = weight_mem_read_arbxbar_arbiters_next_7_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]));
  assign or_556_nl = weight_mem_read_arbxbar_arbiters_next_7_3_sva | nor_tmp_65;
  assign mux_210_nl = MUX_s_1_2_2(or_557_nl, or_556_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign or_555_nl = weight_mem_read_arbxbar_arbiters_next_7_2_sva | or_tmp_225;
  assign mux_211_nl = MUX_s_1_2_2(mux_210_nl, or_555_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign or_554_nl = weight_mem_read_arbxbar_arbiters_next_7_1_sva | and_781_cse
      | or_tmp_225;
  assign mux_tmp_209 = MUX_s_1_2_2(mux_211_nl, or_554_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign or_tmp_232 = and_776_cse | nor_tmp_70;
  assign or_564_nl = Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]));
  assign or_563_nl = Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 | nor_tmp_70;
  assign mux_213_nl = MUX_s_1_2_2(or_564_nl, or_563_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign or_562_nl = Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 | or_tmp_232;
  assign mux_214_nl = MUX_s_1_2_2(mux_213_nl, or_562_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign or_561_nl = Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 | and_777_cse | or_tmp_232;
  assign mux_215_nl = MUX_s_1_2_2(mux_214_nl, or_561_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign mux_216_nl = MUX_s_1_2_2(mux_tmp_209, mux_215_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_558_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7])
      | mux_tmp_209;
  assign mux_217_nl = MUX_s_1_2_2(mux_216_nl, or_558_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_218_nl = MUX_s_1_2_2(mux_tmp_209, mux_217_nl, while_stage_0_5);
  assign and_dcpl_672 = (~ mux_218_nl) & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]))) & nor_285_cse;
  assign and_799_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) & while_mux_1438_tmp;
  assign or_tmp_239 = and_799_cse | (while_mux_1439_tmp & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]));
  assign and_801_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  assign or_tmp_241 = and_801_cse | (weight_mem_read_arbxbar_arbiters_next_6_5_sva
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]));
  assign mux_222_nl = MUX_s_1_2_2(or_tmp_241, or_tmp_239, while_stage_0_5);
  assign or_569_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | or_tmp_241;
  assign or_567_nl = while_mux_1437_tmp | or_tmp_239;
  assign mux_221_nl = MUX_s_1_2_2(or_569_nl, or_567_nl, while_stage_0_5);
  assign mux_tmp_220 = MUX_s_1_2_2(mux_222_nl, mux_221_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign and_805_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & while_mux_1442_tmp;
  assign and_804_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & while_mux_1441_tmp;
  assign and_806_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]) & while_mux_1443_tmp;
  assign nand_10_nl = ~(while_mux_1440_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      & (~ or_tmp_239));
  assign mux_224_nl = MUX_s_1_2_2(nand_10_nl, or_tmp_239, and_804_cse);
  assign mux_225_nl = MUX_s_1_2_2(mux_224_nl, or_tmp_239, and_805_cse);
  assign mux_tmp_223 = MUX_s_1_2_2(mux_225_nl, or_tmp_239, and_806_cse);
  assign and_809_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  assign and_808_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  assign and_810_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  assign nand_11_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      & (~ or_tmp_241));
  assign mux_227_nl = MUX_s_1_2_2(nand_11_nl, or_tmp_241, and_808_cse);
  assign mux_228_nl = MUX_s_1_2_2(mux_227_nl, or_tmp_241, and_809_cse);
  assign mux_tmp_226 = MUX_s_1_2_2(mux_228_nl, or_tmp_241, and_810_cse);
  assign mux_231_nl = MUX_s_1_2_2(mux_tmp_226, mux_tmp_223, while_stage_0_5);
  assign or_571_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | mux_tmp_226;
  assign or_570_nl = while_mux_1437_tmp | mux_tmp_223;
  assign mux_230_nl = MUX_s_1_2_2(or_571_nl, or_570_nl, while_stage_0_5);
  assign mux_232_itm = MUX_s_1_2_2(mux_231_nl, mux_230_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_tmp_246 = ((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]) & while_mux_1437_tmp)
      | and_799_cse;
  assign and_814_cse = while_mux_1440_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign or_576_nl = while_mux_1438_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign or_575_nl = while_mux_1437_tmp | and_799_cse;
  assign mux_233_nl = MUX_s_1_2_2(or_576_nl, or_575_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_234_nl = MUX_s_1_2_2(mux_233_nl, or_tmp_246, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_574_nl = while_mux_1439_tmp | or_tmp_246;
  assign mux_235_nl = MUX_s_1_2_2(mux_234_nl, or_574_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_251 = and_805_cse | and_814_cse | mux_235_nl;
  assign or_tmp_254 = and_801_cse | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  assign mux_tmp_233 = MUX_s_1_2_2(and_801_cse, or_tmp_254, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign and_818_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  assign or_583_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign mux_237_nl = MUX_s_1_2_2(or_583_nl, or_tmp_254, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_238_nl = MUX_s_1_2_2(mux_237_nl, mux_tmp_233, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_582_nl = weight_mem_read_arbxbar_arbiters_next_6_5_sva | mux_tmp_233;
  assign mux_239_nl = MUX_s_1_2_2(mux_238_nl, or_582_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_258 = and_809_cse | and_818_cse | mux_239_nl;
  assign mux_244_nl = MUX_s_1_2_2(or_tmp_258, or_tmp_251, while_stage_0_5);
  assign or_590_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | or_tmp_258;
  assign or_589_nl = while_mux_1441_tmp | or_tmp_251;
  assign mux_243_nl = MUX_s_1_2_2(or_590_nl, or_589_nl, while_stage_0_5);
  assign mux_245_nl = MUX_s_1_2_2(mux_244_nl, mux_243_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign or_588_nl = weight_mem_read_arbxbar_arbiters_next_6_1_sva | or_tmp_258;
  assign or_587_nl = while_mux_1443_tmp | or_tmp_251;
  assign mux_241_nl = MUX_s_1_2_2(or_588_nl, or_587_nl, while_stage_0_5);
  assign or_586_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | or_tmp_258;
  assign or_579_nl = while_mux_1441_tmp | while_mux_1443_tmp | or_tmp_251;
  assign mux_240_nl = MUX_s_1_2_2(or_586_nl, or_579_nl, while_stage_0_5);
  assign mux_242_nl = MUX_s_1_2_2(mux_241_nl, mux_240_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_246_itm = MUX_s_1_2_2(mux_245_nl, mux_242_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_tmp_264 = and_804_cse | and_814_cse;
  assign or_tmp_270 = and_808_cse | and_818_cse;
  assign nor_432_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])));
  assign nor_433_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_3_sva | and_818_cse);
  assign mux_250_nl = MUX_s_1_2_2(nor_432_nl, nor_433_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nor_434_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_2_sva | or_tmp_270);
  assign mux_251_nl = MUX_s_1_2_2(mux_250_nl, nor_434_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign nor_435_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_1_sva | and_809_cse
      | or_tmp_270);
  assign mux_252_nl = MUX_s_1_2_2(mux_251_nl, nor_435_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign nor_436_nl = ~(while_mux_1440_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])));
  assign nor_437_nl = ~(while_mux_1441_tmp | and_814_cse);
  assign mux_247_nl = MUX_s_1_2_2(nor_436_nl, nor_437_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nor_438_nl = ~(while_mux_1442_tmp | or_tmp_264);
  assign mux_248_nl = MUX_s_1_2_2(mux_247_nl, nor_438_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign nor_439_nl = ~(while_mux_1443_tmp | and_805_cse | or_tmp_264);
  assign mux_249_nl = MUX_s_1_2_2(mux_248_nl, nor_439_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign mux_253_nl = MUX_s_1_2_2(mux_252_nl, mux_249_nl, while_stage_0_5);
  assign and_dcpl_675 = mux_253_nl & nor_286_cse & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])));
  assign or_tmp_279 = and_806_cse | and_805_cse | and_804_cse | and_814_cse | or_tmp_239;
  assign or_tmp_284 = and_810_cse | and_809_cse | and_808_cse | and_818_cse | or_tmp_241;
  assign nor_tmp_118 = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]) & while_mux_1432_tmp;
  assign nor_tmp_121 = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  assign and_838_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) & while_mux_1431_tmp;
  assign and_836_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  assign or_614_cse = and_976_cse | and_838_cse | nor_tmp_118;
  assign or_616_cse = and_972_cse | and_836_cse | nor_tmp_121;
  assign mux_tmp_254 = MUX_s_1_2_2(or_616_cse, or_614_cse, while_stage_0_5);
  assign nand_13_nl = ~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_4_sva
      & (~ or_616_cse));
  assign mux_260_itm = MUX_s_1_2_2(nand_13_nl, or_616_cse, and_971_cse);
  assign nand_12_nl = ~(while_mux_1433_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      & (~ or_614_cse));
  assign mux_258_itm = MUX_s_1_2_2(nand_12_nl, or_614_cse, and_975_cse);
  assign mux_270_nl = MUX_s_1_2_2(mux_260_itm, mux_258_itm, while_stage_0_5);
  assign mux_268_nl = MUX_s_1_2_2(mux_260_itm, or_616_cse, weight_mem_read_arbxbar_arbiters_next_5_3_sva);
  assign mux_267_nl = MUX_s_1_2_2(mux_258_itm, or_614_cse, while_mux_1434_tmp);
  assign mux_269_nl = MUX_s_1_2_2(mux_268_nl, mux_267_nl, while_stage_0_5);
  assign mux_271_nl = MUX_s_1_2_2(mux_270_nl, mux_269_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign mux_264_nl = MUX_s_1_2_2(mux_260_itm, or_616_cse, weight_mem_read_arbxbar_arbiters_next_5_1_sva);
  assign mux_263_nl = MUX_s_1_2_2(mux_258_itm, or_614_cse, while_mux_1436_tmp);
  assign mux_265_nl = MUX_s_1_2_2(mux_264_nl, mux_263_nl, while_stage_0_5);
  assign or_620_nl = weight_mem_read_arbxbar_arbiters_next_5_3_sva | weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  assign mux_261_nl = MUX_s_1_2_2(mux_260_itm, or_616_cse, or_620_nl);
  assign or_617_nl = while_mux_1434_tmp | while_mux_1436_tmp;
  assign mux_259_nl = MUX_s_1_2_2(mux_258_itm, or_614_cse, or_617_nl);
  assign mux_262_nl = MUX_s_1_2_2(mux_261_nl, mux_259_nl, while_stage_0_5);
  assign mux_266_nl = MUX_s_1_2_2(mux_265_nl, mux_262_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign mux_272_itm = MUX_s_1_2_2(mux_271_nl, mux_266_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign and_849_cse = while_mux_1436_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign or_tmp_296 = and_849_cse | nor_tmp_118;
  assign or_tmp_297 = and_838_cse | or_tmp_296;
  assign and_851_cse = weight_mem_read_arbxbar_arbiters_next_5_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign or_tmp_304 = and_851_cse | nor_tmp_121;
  assign or_tmp_305 = and_836_cse | or_tmp_304;
  assign mux_276_nl = MUX_s_1_2_2((~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])),
      weight_mem_read_arbxbar_arbiters_next_5_5_sva, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign or_635_nl = and_851_cse | mux_276_nl;
  assign or_634_nl = weight_mem_read_arbxbar_arbiters_next_5_6_sva | or_tmp_304;
  assign mux_277_nl = MUX_s_1_2_2(or_635_nl, or_634_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign or_633_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1
      | or_tmp_305;
  assign mux_278_nl = MUX_s_1_2_2(mux_277_nl, or_633_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign nor_441_nl = ~(and_969_cse | and_970_cse | and_971_cse | mux_278_nl);
  assign mux_273_nl = MUX_s_1_2_2((~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])),
      while_mux_1432_tmp, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign or_627_nl = and_849_cse | mux_273_nl;
  assign or_626_nl = while_mux_1431_tmp | or_tmp_296;
  assign mux_274_nl = MUX_s_1_2_2(or_627_nl, or_626_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign or_625_nl = while_mux_1430_tmp | or_tmp_297;
  assign mux_275_nl = MUX_s_1_2_2(mux_274_nl, or_625_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign nor_442_nl = ~(and_973_cse | and_974_cse | and_975_cse | mux_275_nl);
  assign not_tmp_441 = MUX_s_1_2_2(nor_441_nl, nor_442_nl, while_stage_0_5);
  assign or_tmp_312 = and_975_cse | and_849_cse;
  assign or_tmp_318 = and_971_cse | and_851_cse;
  assign nor_443_nl = ~(weight_mem_read_arbxbar_arbiters_next_5_1_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])));
  assign nor_444_nl = ~(weight_mem_read_arbxbar_arbiters_next_5_2_sva | and_851_cse);
  assign mux_283_nl = MUX_s_1_2_2(nor_443_nl, nor_444_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign nor_445_nl = ~(weight_mem_read_arbxbar_arbiters_next_5_3_sva | or_tmp_318);
  assign mux_284_nl = MUX_s_1_2_2(mux_283_nl, nor_445_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign nor_446_nl = ~(weight_mem_read_arbxbar_arbiters_next_5_4_sva | and_970_cse
      | or_tmp_318);
  assign mux_285_nl = MUX_s_1_2_2(mux_284_nl, nor_446_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign nor_447_nl = ~(while_mux_1436_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])));
  assign nor_448_nl = ~(while_mux_1435_tmp | and_849_cse);
  assign mux_280_nl = MUX_s_1_2_2(nor_447_nl, nor_448_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign nor_449_nl = ~(while_mux_1434_tmp | or_tmp_312);
  assign mux_281_nl = MUX_s_1_2_2(mux_280_nl, nor_449_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign nor_450_nl = ~(while_mux_1433_tmp | and_974_cse | or_tmp_312);
  assign mux_282_nl = MUX_s_1_2_2(mux_281_nl, nor_450_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign mux_286_nl = MUX_s_1_2_2(mux_285_nl, mux_282_nl, while_stage_0_5);
  assign and_dcpl_678 = mux_286_nl & nor_290_cse & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])));
  assign nor_tmp_158 = while_mux_1424_tmp & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign nor_tmp_159 = weight_mem_read_arbxbar_arbiters_next_4_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign or_659_cse = while_mux_1425_tmp | nor_tmp_158;
  assign or_660_cse = weight_mem_read_arbxbar_arbiters_next_4_5_sva | nor_tmp_159;
  assign mux_289_nl = MUX_s_1_2_2(nor_tmp_159, nor_tmp_158, while_stage_0_5);
  assign mux_288_nl = MUX_s_1_2_2(or_660_cse, or_659_cse, while_stage_0_5);
  assign mux_290_nl = MUX_s_1_2_2(mux_289_nl, mux_288_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign or_dcpl_320 = mux_290_nl | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  assign and_869_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]) & while_mux_1427_tmp;
  assign and_870_cse = while_mux_1426_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign or_tmp_335 = and_869_cse | and_870_cse;
  assign and_871_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_1_sva;
  assign and_872_cse = weight_mem_read_arbxbar_arbiters_next_4_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign or_tmp_338 = and_871_cse | and_872_cse | or_tmp_335;
  assign and_874_cse = Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign or_668_nl = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]) & Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1)
      | and_874_cse | or_tmp_335;
  assign mux_292_nl = MUX_s_1_2_2(or_tmp_338, or_668_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign or_664_nl = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4])
      | or_tmp_335;
  assign mux_291_nl = MUX_s_1_2_2(or_tmp_338, or_664_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign mux_tmp_290 = MUX_s_1_2_2(mux_292_nl, mux_291_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_341 = ~((~(while_mux_1424_tmp & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4])))
      & mux_tmp_290);
  assign and_878_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  assign and_879_cse = weight_mem_read_arbxbar_arbiters_next_4_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign or_tmp_345 = and_871_cse | and_872_cse | and_878_cse | and_879_cse;
  assign or_tmp_346 = ~((~(weight_mem_read_arbxbar_arbiters_next_4_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4])))
      & or_tmp_345);
  assign mux_295_nl = MUX_s_1_2_2(or_tmp_346, or_tmp_341, while_stage_0_5);
  assign or_675_nl = weight_mem_read_arbxbar_arbiters_next_4_5_sva | or_tmp_346;
  assign or_670_nl = while_mux_1425_tmp | or_tmp_341;
  assign mux_294_nl = MUX_s_1_2_2(or_675_nl, or_670_nl, while_stage_0_5);
  assign mux_296_nl = MUX_s_1_2_2(mux_295_nl, mux_294_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign and_dcpl_679 = ~(mux_296_nl | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign mux_297_nl = MUX_s_1_2_2(nor_297_cse, while_mux_1424_tmp, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign mux_298_nl = MUX_s_1_2_2(mux_297_nl, or_659_cse, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign or_tmp_352 = and_869_cse | and_870_cse | mux_298_nl;
  assign or_tmp_353 = and_872_cse | or_tmp_352;
  assign or_tmp_355 = and_874_cse | or_tmp_352;
  assign mux_301_nl = MUX_s_1_2_2(nor_297_cse, weight_mem_read_arbxbar_arbiters_next_4_6_sva,
      weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign mux_302_nl = MUX_s_1_2_2(mux_301_nl, or_660_cse, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign or_tmp_361 = and_872_cse | and_878_cse | and_879_cse | mux_302_nl;
  assign mux_304_nl = MUX_s_1_2_2(or_tmp_353, or_tmp_355, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign or_692_nl = (Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_cse
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4])) | or_tmp_352;
  assign mux_305_nl = MUX_s_1_2_2(mux_304_nl, or_692_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_306_nl = MUX_s_1_2_2(or_tmp_361, mux_305_nl, while_stage_0_5);
  assign or_690_nl = weight_mem_read_arbxbar_arbiters_next_4_1_sva | or_tmp_361;
  assign or_685_nl = weight_mem_read_arbxbar_arbiters_next_4_1_sva | or_tmp_353;
  assign or_684_nl = Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 | or_tmp_355;
  assign mux_299_nl = MUX_s_1_2_2(or_685_nl, or_684_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign or_682_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4])
      | weight_mem_read_arbxbar_arbiters_next_4_1_sva | or_tmp_353;
  assign mux_300_nl = MUX_s_1_2_2(mux_299_nl, or_682_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_303_nl = MUX_s_1_2_2(or_690_nl, mux_300_nl, while_stage_0_5);
  assign mux_307_nl = MUX_s_1_2_2(mux_306_nl, mux_303_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign and_dcpl_680 = ~(mux_307_nl | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign or_tmp_369 = and_878_cse | and_879_cse;
  assign or_696_nl = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 | or_tmp_335;
  assign or_695_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4])
      | or_tmp_335;
  assign mux_308_nl = MUX_s_1_2_2(or_696_nl, or_695_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_306 = MUX_s_1_2_2(or_tmp_369, mux_308_nl, while_stage_0_5);
  assign or_700_nl = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4])) | or_tmp_335;
  assign mux_tmp_307 = MUX_s_1_2_2(or_tmp_369, or_700_nl, while_stage_0_5);
  assign or_833_nl = (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1) | or_tmp_335;
  assign mux_311_nl = MUX_s_1_2_2(mux_tmp_307, or_833_nl, weight_mem_read_arbxbar_arbiters_next_4_2_sva);
  assign or_699_nl = weight_mem_read_arbxbar_arbiters_next_4_2_sva | mux_tmp_306;
  assign mux_tmp_309 = MUX_s_1_2_2(mux_311_nl, or_699_nl, Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1);
  assign or_704_nl = weight_mem_read_arbxbar_arbiters_next_4_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]));
  assign or_703_nl = weight_mem_read_arbxbar_arbiters_next_4_3_sva | and_879_cse;
  assign mux_317_nl = MUX_s_1_2_2(or_704_nl, or_703_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign or_702_nl = while_mux_1426_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]));
  assign or_701_nl = while_mux_1427_tmp | and_870_cse;
  assign mux_316_nl = MUX_s_1_2_2(or_702_nl, or_701_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign mux_318_nl = MUX_s_1_2_2(mux_317_nl, mux_316_nl, while_stage_0_5);
  assign mux_319_nl = MUX_s_1_2_2(mux_318_nl, mux_tmp_309, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign mux_313_nl = MUX_s_1_2_2(mux_tmp_307, mux_tmp_309, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign or_698_nl = and_872_cse | mux_tmp_306;
  assign mux_314_nl = MUX_s_1_2_2(mux_313_nl, or_698_nl, Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1);
  assign or_694_nl = Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 | and_874_cse | (~
      while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1) | or_tmp_335;
  assign mux_315_nl = MUX_s_1_2_2(mux_314_nl, or_694_nl, weight_mem_read_arbxbar_arbiters_next_4_1_sva);
  assign mux_320_nl = MUX_s_1_2_2(mux_319_nl, mux_315_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign and_dcpl_684 = ~(mux_320_nl | (~ and_dcpl_593) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]));
  assign or_tmp_377 = nor_tmp_158 | mux_tmp_290;
  assign or_tmp_379 = nor_tmp_159 | or_tmp_345;
  assign and_dcpl_687 = ~(weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp);
  assign nor_tmp_195 = while_mux_1421_tmp & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign or_tmp_381 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]) & while_mux_1422_tmp)
      | nor_tmp_195;
  assign or_tmp_382 = ((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]) & while_mux_1420_tmp)
      | or_tmp_381;
  assign nor_tmp_198 = weight_mem_read_arbxbar_arbiters_next_3_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign or_tmp_384 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_1_sva)
      | nor_tmp_198;
  assign or_tmp_385 = ((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_3_sva)
      | or_tmp_384;
  assign or_716_nl = weight_mem_read_arbxbar_arbiters_next_3_4_sva | or_tmp_385;
  assign Arbiter_8U_Roundrobin_pick_1_mux_610_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1419_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_610_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_713_nl = while_mux_1419_nl | or_tmp_382;
  assign mux_tmp_321 = MUX_s_1_2_2(or_716_nl, or_713_nl, while_stage_0_5);
  assign mux_325_nl = MUX_s_1_2_2(or_tmp_385, or_tmp_382, while_stage_0_5);
  assign mux_tmp_323 = MUX_s_1_2_2(mux_325_nl, mux_tmp_321, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign and_dcpl_688 = mux_tmp_323 & and_dcpl_687;
  assign and_dcpl_689 = (~((~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]))) | mux_tmp_323)) &
      and_dcpl_687;
  assign or_723_nl = weight_mem_read_arbxbar_arbiters_next_3_2_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]));
  assign or_722_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva | nor_tmp_198;
  assign mux_329_nl = MUX_s_1_2_2(or_723_nl, or_722_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign or_721_nl = weight_mem_read_arbxbar_arbiters_next_3_3_sva | or_tmp_384;
  assign mux_330_nl = MUX_s_1_2_2(mux_329_nl, or_721_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign or_720_nl = while_mux_1421_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]));
  assign or_719_nl = while_mux_1422_tmp | nor_tmp_195;
  assign mux_327_nl = MUX_s_1_2_2(or_720_nl, or_719_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign or_718_nl = while_mux_1420_tmp | or_tmp_381;
  assign mux_328_nl = MUX_s_1_2_2(mux_327_nl, or_718_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign mux_331_nl = MUX_s_1_2_2(mux_330_nl, mux_328_nl, while_stage_0_5);
  assign mux_332_nl = MUX_s_1_2_2(mux_331_nl, mux_tmp_321, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign and_dcpl_695 = ~(mux_332_nl | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]));
  assign nor_tmp_200 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  assign and_907_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) & Arbiter_8U_Roundrobin_pick_1_mux_133_mx1w1;
  assign and_909_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_9_mx1w0;
  assign and_908_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) & Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1;
  assign or_725_nl = and_907_cse | and_908_cse;
  assign or_724_nl = and_909_cse | nor_tmp_200;
  assign mux_tmp_330 = MUX_s_1_2_2(or_725_nl, or_724_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_397 = and_736_cse | nor_tmp_200;
  assign mux_335_nl = MUX_s_1_2_2(or_tmp_397, mux_tmp_330, while_stage_0_5);
  assign or_728_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva | or_tmp_397;
  assign or_726_nl = while_mux_1403_tmp | mux_tmp_330;
  assign mux_334_nl = MUX_s_1_2_2(or_728_nl, or_726_nl, while_stage_0_5);
  assign mux_tmp_333 = MUX_s_1_2_2(mux_335_nl, mux_334_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign nor_tmp_209 = while_mux_1406_tmp & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign or_tmp_399 = ((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) & while_mux_1405_tmp)
      | nor_tmp_209;
  assign or_tmp_400 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]) & while_mux_1408_tmp)
      | or_tmp_399;
  assign or_tmp_401 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) & while_mux_1407_tmp)
      | or_tmp_400;
  assign nand_66_cse = ~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1);
  assign or_735_nl = and_907_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      & Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1)) & or_tmp_401));
  assign or_733_nl = and_909_cse | (~(nand_66_cse & or_tmp_401));
  assign mux_tmp_334 = MUX_s_1_2_2(or_735_nl, or_733_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_407 = and_743_cse | and_742_cse;
  assign or_tmp_408 = and_738_cse | or_tmp_407;
  assign or_tmp_409 = and_744_cse | or_tmp_408;
  assign or_tmp_411 = and_736_cse | (~(nand_66_cse & or_tmp_409));
  assign mux_339_nl = MUX_s_1_2_2(or_tmp_411, mux_tmp_334, while_stage_0_5);
  assign or_742_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva | or_tmp_411;
  assign or_736_nl = while_mux_1403_tmp | mux_tmp_334;
  assign mux_338_nl = MUX_s_1_2_2(or_742_nl, or_736_nl, while_stage_0_5);
  assign mux_340_itm = MUX_s_1_2_2(mux_339_nl, mux_338_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign or_tmp_413 = nor_tmp_200 | or_tmp_401;
  assign or_tmp_415 = and_908_cse | or_tmp_401;
  assign or_746_nl = and_907_cse | or_tmp_415;
  assign or_744_nl = and_909_cse | or_tmp_413;
  assign mux_tmp_338 = MUX_s_1_2_2(or_746_nl, or_744_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_418 = nor_tmp_200 | or_tmp_409;
  assign or_tmp_419 = and_736_cse | or_tmp_418;
  assign or_750_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva | or_tmp_419;
  assign or_747_nl = while_mux_1403_tmp | mux_tmp_338;
  assign mux_tmp_339 = MUX_s_1_2_2(or_750_nl, or_747_nl, while_stage_0_5);
  assign nand_tmp_17 = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) & (~
      or_tmp_401));
  assign nand_18_nl = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) & (~
      or_tmp_409));
  assign or_756_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      | or_tmp_409;
  assign mux_348_nl = MUX_s_1_2_2(nand_18_nl, or_756_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign or_755_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_418;
  assign mux_349_nl = MUX_s_1_2_2(mux_348_nl, or_755_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign or_754_nl = Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 | or_tmp_401;
  assign mux_345_nl = MUX_s_1_2_2(nand_tmp_17, or_754_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign or_753_nl = Arbiter_8U_Roundrobin_pick_1_mux_133_mx1w1 | or_tmp_415;
  assign mux_346_nl = MUX_s_1_2_2(mux_345_nl, or_753_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign or_752_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      | or_tmp_401;
  assign mux_343_nl = MUX_s_1_2_2(nand_tmp_17, or_752_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign or_751_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_9_mx1w0
      | or_tmp_413;
  assign mux_344_nl = MUX_s_1_2_2(mux_343_nl, or_751_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign mux_347_nl = MUX_s_1_2_2(mux_346_nl, mux_344_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_350_nl = MUX_s_1_2_2(mux_349_nl, mux_347_nl, while_stage_0_5);
  assign mux_351_itm = MUX_s_1_2_2(mux_350_nl, mux_tmp_339, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign nor_463_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_3_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])));
  assign nor_464_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_4_sva | and_742_cse);
  assign mux_355_nl = MUX_s_1_2_2(nor_463_nl, nor_464_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign nor_465_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_1_sva | or_tmp_407);
  assign mux_356_nl = MUX_s_1_2_2(mux_355_nl, nor_465_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign nor_466_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_2_sva | or_tmp_408);
  assign mux_357_nl = MUX_s_1_2_2(mux_356_nl, nor_466_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign nor_467_nl = ~(while_mux_1406_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])));
  assign nor_468_nl = ~(while_mux_1405_tmp | nor_tmp_209);
  assign mux_352_nl = MUX_s_1_2_2(nor_467_nl, nor_468_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign nor_469_nl = ~(while_mux_1408_tmp | or_tmp_399);
  assign mux_353_nl = MUX_s_1_2_2(mux_352_nl, nor_469_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign nor_470_nl = ~(while_mux_1407_tmp | or_tmp_400);
  assign mux_354_nl = MUX_s_1_2_2(mux_353_nl, nor_470_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign mux_358_nl = MUX_s_1_2_2(mux_357_nl, mux_354_nl, while_stage_0_5);
  assign and_dcpl_697 = mux_358_nl & and_dcpl_615;
  assign nor_tmp_224 = while_mux_1396_tmp & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign or_tmp_436 = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0])
      | weight_mem_read_arbxbar_arbiters_next_0_5_sva | nor_tmp_224;
  assign mux_tmp_358 = MUX_s_1_2_2(nor_tmp_224, or_tmp_436, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign or_769_nl = weight_mem_read_arbxbar_arbiters_next_0_5_sva | nor_tmp_224;
  assign or_768_nl = Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 | nor_tmp_224;
  assign mux_tmp_359 = MUX_s_1_2_2(or_769_nl, or_768_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign mux_tmp_360 = MUX_s_1_2_2(nor_tmp_224, mux_tmp_359, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign mux_365_nl = MUX_s_1_2_2(mux_tmp_360, mux_tmp_358, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_770_nl = Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 | mux_tmp_360;
  assign or_767_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | mux_tmp_358;
  assign mux_364_nl = MUX_s_1_2_2(or_770_nl, or_767_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_363 = MUX_s_1_2_2(mux_365_nl, mux_364_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign nor_tmp_227 = weight_mem_read_arbxbar_arbiters_next_0_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign or_tmp_441 = ((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) & weight_mem_read_arbxbar_arbiters_next_0_5_sva)
      | nor_tmp_227;
  assign or_tmp_442 = and_979_cse | or_tmp_441;
  assign mux_tmp_364 = MUX_s_1_2_2(or_tmp_442, mux_tmp_363, while_stage_0_5);
  assign and_936_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]) & while_mux_1401_tmp;
  assign nand_19_nl = ~(while_mux_1400_tmp & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0])
      & (~ mux_tmp_358));
  assign mux_tmp_365 = MUX_s_1_2_2(nand_19_nl, mux_tmp_358, and_936_cse);
  assign nand_20_nl = ~(while_mux_1400_tmp & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0])
      & (~ mux_tmp_360));
  assign mux_tmp_366 = MUX_s_1_2_2(nand_20_nl, mux_tmp_360, and_936_cse);
  assign and_941_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]) & weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  assign nand_21_nl = ~(weight_mem_read_arbxbar_arbiters_next_0_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0])
      & (~ or_tmp_441));
  assign mux_375_nl = MUX_s_1_2_2(nand_21_nl, or_tmp_441, and_941_cse);
  assign or_775_nl = and_979_cse | mux_375_nl;
  assign mux_376_nl = MUX_s_1_2_2(or_775_nl, or_tmp_442, and_978_cse);
  assign mux_377_nl = MUX_s_1_2_2(mux_376_nl, or_tmp_442, and_977_cse);
  assign mux_371_nl = MUX_s_1_2_2(mux_tmp_366, mux_tmp_365, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_774_nl = Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 | mux_tmp_366;
  assign or_773_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | mux_tmp_365;
  assign mux_370_nl = MUX_s_1_2_2(or_774_nl, or_773_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_372_nl = MUX_s_1_2_2(mux_371_nl, mux_370_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign mux_373_nl = MUX_s_1_2_2(mux_372_nl, mux_tmp_363, and_981_cse);
  assign mux_374_nl = MUX_s_1_2_2(mux_373_nl, mux_tmp_363, and_980_cse);
  assign mux_378_itm = MUX_s_1_2_2(mux_377_nl, mux_374_nl, while_stage_0_5);
  assign and_947_cse = while_mux_1400_tmp & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign or_tmp_447 = and_936_cse | and_947_cse | mux_tmp_358;
  assign or_tmp_450 = and_936_cse | and_947_cse | mux_tmp_360;
  assign or_781_nl = Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 | or_tmp_450;
  assign or_778_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | or_tmp_447;
  assign mux_tmp_376 = MUX_s_1_2_2(or_781_nl, or_778_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_452 = (~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])) |
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign mux_tmp_377 = MUX_s_1_2_2(nor_310_cse, or_tmp_452, while_mux_1396_tmp);
  assign and_951_cse = weight_mem_read_arbxbar_arbiters_next_0_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign or_tmp_460 = and_941_cse | and_951_cse | or_tmp_441;
  assign mux_385_nl = MUX_s_1_2_2(nor_310_cse, or_tmp_452, weight_mem_read_arbxbar_arbiters_next_0_6_sva);
  assign or_792_nl = weight_mem_read_arbxbar_arbiters_next_0_5_sva | nor_tmp_227;
  assign mux_386_nl = MUX_s_1_2_2(mux_385_nl, or_792_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign or_794_nl = and_941_cse | and_951_cse | mux_386_nl;
  assign or_791_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | or_tmp_460;
  assign mux_387_nl = MUX_s_1_2_2(or_794_nl, or_791_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign nor_471_nl = ~(and_977_cse | and_978_cse | mux_387_nl);
  assign mux_382_nl = MUX_s_1_2_2(mux_tmp_377, mux_tmp_359, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign or_786_nl = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]) & Arbiter_8U_Roundrobin_pick_1_mux_63_mx1w1)
      | (Arbiter_8U_Roundrobin_pick_1_mux_62_mx1w1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]))
      | mux_382_nl;
  assign mux_381_nl = MUX_s_1_2_2(mux_tmp_377, or_tmp_436, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign or_784_nl = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0)
      | (Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]))
      | mux_381_nl;
  assign mux_383_nl = MUX_s_1_2_2(or_786_nl, or_784_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_384_nl = MUX_s_1_2_2(mux_383_nl, mux_tmp_376, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign nor_472_nl = ~(and_980_cse | and_981_cse | mux_384_nl);
  assign not_tmp_470 = MUX_s_1_2_2(nor_471_nl, nor_472_nl, while_stage_0_5);
  assign or_tmp_467 = and_936_cse | and_947_cse;
  assign or_tmp_473 = and_941_cse | and_951_cse;
  assign nor_473_nl = ~(weight_mem_read_arbxbar_arbiters_next_0_2_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0])));
  assign nor_474_nl = ~(weight_mem_read_arbxbar_arbiters_next_0_1_sva | and_951_cse);
  assign mux_392_nl = MUX_s_1_2_2(nor_473_nl, nor_474_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]);
  assign nor_475_nl = ~(weight_mem_read_arbxbar_arbiters_next_0_3_sva | or_tmp_473);
  assign mux_393_nl = MUX_s_1_2_2(mux_392_nl, nor_475_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign nor_476_nl = ~(weight_mem_read_arbxbar_arbiters_next_0_4_sva | and_978_cse
      | or_tmp_473);
  assign mux_394_nl = MUX_s_1_2_2(mux_393_nl, nor_476_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign nor_477_nl = ~(while_mux_1400_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0])));
  assign nor_478_nl = ~(while_mux_1401_tmp | and_947_cse);
  assign mux_389_nl = MUX_s_1_2_2(nor_477_nl, nor_478_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]);
  assign nor_479_nl = ~(while_mux_1399_tmp | or_tmp_467);
  assign mux_390_nl = MUX_s_1_2_2(mux_389_nl, nor_479_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign nor_480_nl = ~(while_mux_1398_tmp | and_981_cse | or_tmp_467);
  assign mux_391_nl = MUX_s_1_2_2(mux_390_nl, nor_480_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign mux_395_nl = MUX_s_1_2_2(mux_394_nl, mux_391_nl, while_stage_0_5);
  assign and_dcpl_700 = mux_395_nl & nor_310_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])));
  assign and_dcpl_704 = (~(weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp))
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp)
      & weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp;
  assign and_dcpl_705 = ~((~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]))) | weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_dcpl_708 = nor_302_cse & (~ (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]))
      & (~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]) | weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp));
  assign or_dcpl_328 = ~(Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs);
  assign ProductSum_for_acc_20_cmp_a = weight_port_read_out_data_7_1_sva_dfm_2;
  assign ProductSum_for_acc_20_cmp_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[15:8];
  assign ProductSum_for_acc_20_cmp_load = ProductSum_for_asn_28_itm_5;
  assign ProductSum_for_acc_20_cmp_datavalid_pff = and_dcpl_35;
  assign ProductSum_for_acc_19_cmp_a0 = weight_port_read_out_data_7_2_sva_dfm_1;
  assign ProductSum_for_acc_19_cmp_a1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[23:16];
  assign ProductSum_for_acc_19_cmp_b0 = weight_port_read_out_data_7_3_sva_dfm_1;
  assign ProductSum_for_acc_19_cmp_b1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[31:24];
  assign ProductSum_for_acc_19_cmp_c0 = weight_port_read_out_data_7_0_sva_dfm_1;
  assign ProductSum_for_acc_19_cmp_c1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[7:0];
  assign ProductSum_for_acc_19_cmp_load_pff = ProductSum_for_asn_26_itm_6;
  assign ProductSum_for_acc_19_cmp_datavalid_pff = and_dcpl_507;
  assign ProductSum_for_acc_18_cmp_a0 = weight_port_read_out_data_7_7_sva_dfm_1;
  assign ProductSum_for_acc_18_cmp_a1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[63:56];
  assign ProductSum_for_acc_18_cmp_b0 = weight_port_read_out_data_7_4_sva_dfm_1;
  assign ProductSum_for_acc_18_cmp_b1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[39:32];
  assign ProductSum_for_acc_18_cmp_c0 = weight_port_read_out_data_7_5_sva_dfm_1;
  assign ProductSum_for_acc_18_cmp_c1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[47:40];
  assign ProductSum_for_acc_17_cmp_a0 = weight_port_read_out_data_7_8_sva_dfm_1;
  assign ProductSum_for_acc_17_cmp_a1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[71:64];
  assign ProductSum_for_acc_17_cmp_b0 = weight_port_read_out_data_7_9_sva_dfm_1;
  assign ProductSum_for_acc_17_cmp_b1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[79:72];
  assign ProductSum_for_acc_17_cmp_c0 = weight_port_read_out_data_7_6_sva_dfm_1;
  assign ProductSum_for_acc_17_cmp_c1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[55:48];
  assign ProductSum_for_acc_16_cmp_a0 = weight_port_read_out_data_7_13_sva_dfm_1;
  assign ProductSum_for_acc_16_cmp_a1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[111:104];
  assign ProductSum_for_acc_16_cmp_b0 = weight_port_read_out_data_7_10_sva_dfm_1;
  assign ProductSum_for_acc_16_cmp_b1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[87:80];
  assign ProductSum_for_acc_16_cmp_c0 = weight_port_read_out_data_7_11_sva_dfm_1;
  assign ProductSum_for_acc_16_cmp_c1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[95:88];
  assign ProductSum_for_acc_15_cmp_a0 = weight_port_read_out_data_7_14_sva_dfm_1;
  assign ProductSum_for_acc_15_cmp_a1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[119:112];
  assign ProductSum_for_acc_15_cmp_b0 = weight_port_read_out_data_7_15_sva_dfm_1;
  assign ProductSum_for_acc_15_cmp_b1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[127:120];
  assign ProductSum_for_acc_15_cmp_c0 = weight_port_read_out_data_7_12_sva_dfm_1;
  assign ProductSum_for_acc_15_cmp_c1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[103:96];
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_6_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_load = ProductSum_for_asn_41_itm_5;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_a0 = weight_mem_run_3_for_5_mux_98_itm_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_b0 = weight_mem_run_3_for_5_mux_99_itm_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_c0 = weight_mem_run_3_for_5_mux_96_itm_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_pff = ProductSum_for_asn_40_itm_6;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a0 = rva_out_reg_data_71_64_sva_dfm_4_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_b0 = {rva_out_reg_data_111_104_sva_dfm_4_1_7
      , rva_out_reg_data_111_104_sva_dfm_4_1_6_0};
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_c0 = {rva_out_reg_data_119_112_sva_dfm_4_1_7
      , rva_out_reg_data_119_112_sva_dfm_4_1_6_0};
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a0 = rva_out_reg_data_79_72_sva_dfm_4_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_b0 = {rva_out_reg_data_87_80_sva_dfm_4_1_7_4
      , rva_out_reg_data_87_80_sva_dfm_4_1_3_0};
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_c0 = {rva_out_reg_data_127_120_sva_dfm_4_1_7_6
      , rva_out_reg_data_127_120_sva_dfm_4_1_5_0};
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0 = {weight_mem_run_3_for_5_mux_109_itm_1_7_6
      , weight_mem_run_3_for_5_mux_109_itm_1_5_0};
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0 = rva_out_reg_data_95_88_sva_dfm_4_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0 = {weight_mem_run_3_for_5_mux_107_itm_1_7
      , weight_mem_run_3_for_5_mux_107_itm_1_6_0};
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0 = {weight_mem_run_3_for_5_mux_110_itm_1_7
      , weight_mem_run_3_for_5_mux_110_itm_1_6_0};
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0 = {weight_mem_run_3_for_5_mux_111_itm_1_7
      , weight_mem_run_3_for_5_mux_111_itm_1_6_0};
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0 = {weight_mem_run_3_for_5_mux_108_itm_1_7
      , weight_mem_run_3_for_5_mux_108_itm_1_6_0};
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_5_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_load = ProductSum_for_asn_56_itm_5;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_a0 = weight_mem_run_3_for_5_mux_82_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_b0 = weight_mem_run_3_for_5_mux_83_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_c0 = weight_mem_run_3_for_5_mux_80_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_pff = ProductSum_for_asn_55_itm_6;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a0 = weight_mem_run_3_for_5_mux_87_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_b0 = weight_mem_run_3_for_5_mux_84_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_c0 = weight_mem_run_3_for_5_mux_85_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a0 = weight_mem_run_3_for_5_mux_88_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_b0 = weight_mem_run_3_for_5_mux_89_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_c0 = weight_mem_run_3_for_5_mux_86_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0 = weight_mem_run_3_for_5_mux_93_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0 = weight_mem_run_3_for_5_mux_90_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0 = weight_mem_run_3_for_5_mux_91_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0 = weight_port_read_out_data_5_14_sva_dfm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0 = weight_port_read_out_data_5_15_sva_dfm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0 = weight_mem_run_3_for_5_mux_92_itm_1;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_port_read_out_data_4_1_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[15:8];
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_pff = ProductSum_for_asn_69_itm_6;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
      weight_port_read_out_data_4_2_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
      weight_port_read_out_data_4_3_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
      weight_port_read_out_data_4_0_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
      weight_port_read_out_data_4_7_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
      weight_port_read_out_data_4_4_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
      weight_port_read_out_data_4_5_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
      weight_port_read_out_data_4_8_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
      weight_port_read_out_data_4_9_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
      weight_port_read_out_data_4_6_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
      weight_port_read_out_data_4_13_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
      weight_port_read_out_data_4_10_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
      weight_port_read_out_data_4_11_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
      weight_port_read_out_data_4_14_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0 = weight_mem_run_3_for_5_mux_79_itm_1;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014,
      weight_port_read_out_data_4_12_sva_dfm_1, and_dcpl_541);
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_3_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_load = ProductSum_for_asn_82_itm_5;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_a0 = weight_mem_run_3_for_5_mux_50_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_b0 = weight_mem_run_3_for_5_mux_51_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_c0 = weight_mem_run_3_for_5_mux_48_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_pff = ProductSum_for_asn_81_itm_6;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a0 = weight_mem_run_3_for_5_mux_55_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_b0 = weight_mem_run_3_for_5_mux_52_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_c0 = weight_mem_run_3_for_5_mux_53_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a0 = weight_mem_run_3_for_5_mux_56_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_b0 = weight_mem_run_3_for_5_mux_57_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_c0 = weight_mem_run_3_for_5_mux_54_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0 = weight_mem_run_3_for_5_mux_61_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0 = weight_mem_run_3_for_5_mux_58_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0 = weight_mem_run_3_for_5_mux_59_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0 = weight_mem_run_3_for_5_mux_62_itm_1;
  assign and_552_nl = fsm_output & (~ weight_mem_run_3_for_land_4_lpi_1_dfm_3);
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000,
      weight_port_read_out_data_3_15_sva_dfm_1, and_552_nl);
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0 = weight_mem_run_3_for_5_mux_60_itm_1;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_port_read_out_data_2_1_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_pff = ProductSum_for_asn_95_itm_6;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
      weight_port_read_out_data_2_2_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
      weight_port_read_out_data_2_3_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
      weight_port_read_out_data_2_0_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
      weight_port_read_out_data_2_7_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
      weight_port_read_out_data_2_4_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
      weight_port_read_out_data_2_5_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
      weight_port_read_out_data_2_8_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
      weight_port_read_out_data_2_9_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
      weight_port_read_out_data_2_6_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
      weight_port_read_out_data_2_13_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
      weight_port_read_out_data_2_10_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
      weight_port_read_out_data_2_11_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
      weight_port_read_out_data_2_14_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0 = weight_mem_run_3_for_5_mux_47_itm_1;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014,
      weight_port_read_out_data_2_12_sva_dfm_1, and_dcpl_539);
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_1_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_load = ProductSum_for_asn_108_itm_5;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_a0 = weight_mem_run_3_for_5_mux_18_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_b0 = weight_mem_run_3_for_5_mux_19_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_c0 = weight_mem_run_3_for_5_mux_16_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_pff = ProductSum_for_asn_107_itm_6;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a0 = weight_mem_run_3_for_5_mux_23_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_b0 = weight_mem_run_3_for_5_mux_20_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_c0 = weight_mem_run_3_for_5_mux_21_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a0 = weight_mem_run_3_for_5_mux_24_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_b0 = weight_mem_run_3_for_5_mux_25_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_c0 = weight_mem_run_3_for_5_mux_22_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0 = weight_mem_run_3_for_5_mux_29_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0 = weight_mem_run_3_for_5_mux_26_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0 = weight_mem_run_3_for_5_mux_27_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0 = weight_mem_run_3_for_5_mux_30_itm_1;
  assign and_550_nl = fsm_output & (~ weight_mem_run_3_for_land_2_lpi_1_dfm_3);
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0 = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000,
      weight_port_read_out_data_1_15_sva_dfm_1, and_550_nl);
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0 = weight_mem_run_3_for_5_mux_28_itm_1;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_a = MUX_v_8_2_2(({weight_port_read_out_data_0_1_sva_mx0_7_4
      , weight_port_read_out_data_0_1_sva_mx0_3_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_load = ProductSum_for_asn_128_itm_5;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_a0 = {weight_port_read_out_data_0_2_sva_dfm_1_1_7
      , weight_port_read_out_data_0_2_sva_dfm_1_1_6_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_b0 = {weight_port_read_out_data_0_3_sva_dfm_1_1_7
      , weight_port_read_out_data_0_3_sva_dfm_1_1_6_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_c0 = {weight_port_read_out_data_0_0_sva_dfm_1_1_7_4
      , weight_port_read_out_data_0_0_sva_dfm_1_1_3_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_pff = ProductSum_for_asn_126_itm_6;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a0 = weight_port_read_out_data_0_7_sva_dfm_1_1;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_b0 = {weight_port_read_out_data_0_4_sva_dfm_1_1_7_4
      , weight_port_read_out_data_0_4_sva_dfm_1_1_3_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_c0 = weight_port_read_out_data_0_5_sva_dfm_1_1;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a0 = weight_mem_run_3_for_5_mux_8_itm_1;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_b0 = weight_mem_run_3_for_5_mux_9_itm_1;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_c0 = weight_mem_run_3_for_5_mux_6_itm_1;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0 = {weight_mem_run_3_for_5_mux_13_itm_1_7
      , weight_mem_run_3_for_5_mux_13_itm_1_6_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0 = {rva_out_reg_data_103_96_sva_dfm_4_1_7_4
      , rva_out_reg_data_103_96_sva_dfm_4_1_3_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0 = {weight_mem_run_3_for_5_mux_11_itm_1_7
      , weight_mem_run_3_for_5_mux_11_itm_1_6_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0 = {weight_mem_run_3_for_5_mux_14_itm_1_7
      , weight_mem_run_3_for_5_mux_14_itm_1_6_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0 = {weight_mem_run_3_for_5_mux_15_itm_1_7_6
      , weight_mem_run_3_for_5_mux_15_itm_1_5_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0 = {weight_mem_run_3_for_5_mux_12_itm_1_7_6
      , weight_mem_run_3_for_5_mux_12_itm_1_5_0};
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0));
  assign weight_mem_banks_write_if_for_if_and_35_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_36_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_37_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_38_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_39_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_40_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_41_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      , weight_mem_banks_write_if_for_if_and_35_nl , weight_mem_banks_write_if_for_if_and_36_nl
      , weight_mem_banks_write_if_for_if_and_37_nl , weight_mem_banks_write_if_for_if_and_38_nl
      , weight_mem_banks_write_if_for_if_and_39_nl , weight_mem_banks_write_if_for_if_and_40_nl
      , weight_mem_banks_write_if_for_if_and_41_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0});
  assign weight_mem_banks_write_if_for_if_mux_7_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      , weight_mem_banks_write_if_for_if_mux_7_nl};
  assign nor_497_nl = ~((~ PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3) |
      PECore_RunFSM_switch_lp_equal_tmp_1_2);
  assign mux_146_nl = MUX_s_1_2_2(mux_tmp_118, nor_497_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff = mux_146_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_2[14:3];
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff = and_dcpl_171;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0));
  assign weight_mem_banks_write_if_for_if_and_28_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_29_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_30_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_31_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_32_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_33_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_34_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      , weight_mem_banks_write_if_for_if_and_28_nl , weight_mem_banks_write_if_for_if_and_29_nl
      , weight_mem_banks_write_if_for_if_and_30_nl , weight_mem_banks_write_if_for_if_and_31_nl
      , weight_mem_banks_write_if_for_if_and_32_nl , weight_mem_banks_write_if_for_if_and_33_nl
      , weight_mem_banks_write_if_for_if_and_34_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0});
  assign weight_mem_banks_write_if_for_if_mux_6_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      , weight_mem_banks_write_if_for_if_mux_6_nl};
  assign nor_496_nl = ~((~ PECore_RunMac_PECore_RunMac_if_and_svs_3) | PECore_UpdateFSM_switch_lp_equal_tmp_2_3);
  assign mux_145_nl = MUX_s_1_2_2(or_85_cse, nor_496_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff = mux_145_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff = and_dcpl_175;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0));
  assign weight_mem_banks_write_if_for_if_and_21_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_22_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_23_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_24_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_25_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_26_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_27_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      , weight_mem_banks_write_if_for_if_and_21_nl , weight_mem_banks_write_if_for_if_and_22_nl
      , weight_mem_banks_write_if_for_if_and_23_nl , weight_mem_banks_write_if_for_if_and_24_nl
      , weight_mem_banks_write_if_for_if_and_25_nl , weight_mem_banks_write_if_for_if_and_26_nl
      , weight_mem_banks_write_if_for_if_and_27_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0});
  assign weight_mem_banks_write_if_for_if_mux_5_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      , weight_mem_banks_write_if_for_if_mux_5_nl};
  assign nor_495_nl = ~((~ PECore_RunMac_PECore_RunMac_if_and_svs_st_3) | ProductSum_for_asn_108_itm_3);
  assign mux_144_nl = MUX_s_1_2_2(or_92_cse, nor_495_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff = mux_144_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff = and_dcpl_178;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0));
  assign weight_mem_banks_write_if_for_if_and_14_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_15_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_16_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_17_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_18_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_19_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_20_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      , weight_mem_banks_write_if_for_if_and_14_nl , weight_mem_banks_write_if_for_if_and_15_nl
      , weight_mem_banks_write_if_for_if_and_16_nl , weight_mem_banks_write_if_for_if_and_17_nl
      , weight_mem_banks_write_if_for_if_and_18_nl , weight_mem_banks_write_if_for_if_and_19_nl
      , weight_mem_banks_write_if_for_if_and_20_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0});
  assign weight_mem_banks_write_if_for_if_mux_4_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      , weight_mem_banks_write_if_for_if_mux_4_nl};
  assign nor_494_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_3) | ProductSum_for_asn_128_itm_3);
  assign mux_143_nl = MUX_s_1_2_2(mux_tmp_108, nor_494_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff = mux_143_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff = and_dcpl_182;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0));
  assign weight_mem_banks_write_if_for_if_and_7_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_9_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_10_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_11_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_12_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_13_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      , weight_mem_banks_write_if_for_if_and_7_nl , weight_mem_banks_write_if_for_if_and_8_nl
      , weight_mem_banks_write_if_for_if_and_9_nl , weight_mem_banks_write_if_for_if_and_10_nl
      , weight_mem_banks_write_if_for_if_and_11_nl , weight_mem_banks_write_if_for_if_and_12_nl
      , weight_mem_banks_write_if_for_if_and_13_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0});
  assign weight_mem_banks_write_if_for_if_mux_3_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      , weight_mem_banks_write_if_for_if_mux_3_nl};
  assign nor_493_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3) | ProductSum_for_asn_28_itm_3);
  assign mux_142_nl = MUX_s_1_2_2(or_106_cse, nor_493_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff = mux_142_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff = and_dcpl_187;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0));
  assign weight_mem_banks_write_if_for_if_and_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_1_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_2_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_3_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_5_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl ,
      weight_mem_banks_write_if_for_if_and_nl , weight_mem_banks_write_if_for_if_and_1_nl
      , weight_mem_banks_write_if_for_if_and_2_nl , weight_mem_banks_write_if_for_if_and_3_nl
      , weight_mem_banks_write_if_for_if_and_4_nl , weight_mem_banks_write_if_for_if_and_5_nl
      , weight_mem_banks_write_if_for_if_and_6_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0});
  assign weight_mem_banks_write_if_for_if_mux_2_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      , weight_mem_banks_write_if_for_if_mux_2_nl};
  assign nor_492_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1)
      | ProductSum_for_asn_41_itm_3);
  assign mux_141_nl = MUX_s_1_2_2(or_113_cse, nor_492_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff = mux_141_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff = and_dcpl_191;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_14_lpi_1_dfm_1_3_2 , weight_write_data_data_0_13_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_12_lpi_1_dfm_1_3_2 , weight_write_data_data_0_11_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_10_lpi_1_dfm_1_3_2 , weight_write_data_data_0_9_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_8_lpi_1_dfm_1_3_2 , weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_1_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_54_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0,
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_1_nl
      , weight_mem_banks_write_if_for_if_mux_54_nl};
  assign nor_491_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1);
  assign mux_140_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_491_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff = mux_140_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_3_14_3;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff = and_dcpl_516;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_14_lpi_1_dfm_1_3_2 , weight_write_data_data_0_13_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_12_lpi_1_dfm_1_3_2 , weight_write_data_data_0_11_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_10_lpi_1_dfm_1_3_2 , weight_write_data_data_0_9_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_8_lpi_1_dfm_1_3_2 , weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_53_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0,
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_nl
      , weight_mem_banks_write_if_for_if_mux_53_nl};
  assign nor_490_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1);
  assign mux_139_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_490_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff = mux_139_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff = and_dcpl_514;
  assign and_dcpl = (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1;
  assign and_dcpl_709 = (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1;
  assign or_dcpl = and_dcpl_709 | and_dcpl;
  assign or_dcpl_329 = and_dcpl_709 | ((pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1);
  assign or_dcpl_331 = ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]) & and_dcpl_634)
      | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]) & and_dcpl_633) | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1])
      & and_dcpl_631);
  assign or_dcpl_333 = ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]) & and_dcpl_638)
      | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]) & and_dcpl_637) | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1])
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]));
  assign or_dcpl_334 = ((~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1])) &
      (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]) & nor_tmp_2)
      | (nor_352_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign and_dcpl_721 = or_dcpl_333 & nor_tmp_2;
  assign and_651_ssc = nor_tmp_2 & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign and_652_ssc = nor_tmp_2 & and_dcpl_637;
  assign and_653_ssc = nor_tmp_2 & and_dcpl_638;
  assign and_655_ssc = (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      & weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_658_ssc = nor_352_cse & (~(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4));
  assign and_661_ssc = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign PECore_DecodeAxiRead_switch_lp_mux_23_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[0]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl
      = PECore_DecodeAxiRead_switch_lp_mux_23_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_37_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl,
      rva_out_reg_data_0_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_24_itm = MUX_s_1_2_2(rva_out_reg_data_mux_37_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_DecodeAxiRead_switch_lp_mux_24_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[8]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl
      = PECore_DecodeAxiRead_switch_lp_mux_24_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_38_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl,
      rva_out_reg_data_8_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_25_itm = MUX_s_1_2_2(rva_out_reg_data_mux_38_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_DecodeAxiRead_switch_lp_mux_25_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[16]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl
      = PECore_DecodeAxiRead_switch_lp_mux_25_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_39_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl,
      rva_out_reg_data_16_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_26_itm = MUX_s_1_2_2(rva_out_reg_data_mux_39_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_DecodeAxiRead_switch_lp_mux_26_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[24]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl
      = PECore_DecodeAxiRead_switch_lp_mux_26_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_41_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl,
      rva_out_reg_data_24_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_27_nl = MUX_s_1_2_2(rva_out_reg_data_mux_41_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_PushAxiRsp_if_mux1h_15 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_27_nl,
      (weight_port_read_out_data_0_3_sva_dfm_4_6_0[0]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign PECore_DecodeAxiRead_switch_lp_mux_22_nl = MUX_v_6_2_2((SC_SRAM_CONFIG[30:25]),
      rva_out_reg_data_30_25_sva_dfm_7, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl =
      MUX_v_6_2_2(6'b000000, PECore_DecodeAxiRead_switch_lp_mux_22_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_16 = MUX1HOT_v_6_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl,
      rva_out_reg_data_30_25_sva_dfm_6, input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4,
      (weight_port_read_out_data_0_3_sva_dfm_4_6_0[6:1]), {PECore_PushAxiRsp_if_asn_79
      , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl
      = (SC_SRAM_CONFIG[31]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8) &
      PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_40_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl,
      rva_out_reg_data_31_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_28_nl = MUX_s_1_2_2(rva_out_reg_data_mux_40_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_PushAxiRsp_if_mux1h_17 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_28_nl,
      weight_port_read_out_data_0_3_sva_dfm_4_7, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign mux_10_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_5, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_11_nl = MUX_s_1_2_2(mux_10_nl, (~ or_tmp_15), or_tmp_14);
  assign weight_mem_run_3_for_5_and_199_ssc = PECoreRun_wen & mux_11_nl & while_stage_0_7;
  assign nor_279_nl = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      | rva_in_reg_rw_sva_st_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5
      | (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4) | PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      | rva_in_reg_rw_sva_5);
  assign mux_12_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_5, nor_279_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_13_nl = MUX_s_1_2_2(mux_12_nl, (~ or_tmp_15), or_tmp_14);
  assign weight_mem_run_3_for_5_and_202_ssc = PECoreRun_wen & mux_13_nl & while_stage_0_7;
  assign weight_port_read_out_data_and_136_ssc = PECoreRun_wen & (~(mux_15_itm &
      (~((~ rva_in_reg_rw_sva_st_1_5) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3))
      & while_stage_0_6)) & and_dcpl_47;
  assign and_1607_cse = weight_mem_run_3_for_land_1_lpi_1_dfm_2 & while_stage_0_6;
  assign and_1608_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & while_stage_0_6;
  assign mux_524_nl = MUX_s_1_2_2((~ mux_522_cse), or_tmp_584, and_1607_cse);
  assign mux_523_nl = MUX_s_1_2_2((~ mux_522_cse), or_tmp_584, and_1608_cse);
  assign mux_525_nl = MUX_s_1_2_2(mux_524_nl, mux_523_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_1529_cse = (~ mux_525_nl) & and_dcpl_47 & PECoreRun_wen;
  assign and_1022_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_dcpl_329);
  assign mux_31_nl = MUX_s_1_2_2(or_tmp_23, (~ or_tmp_37), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_30_nl = MUX_s_1_2_2((~ or_tmp_37), or_tmp_23, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_32_nl = MUX_s_1_2_2(mux_31_nl, mux_30_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign or_191_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])
      | (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_29_nl = MUX_s_1_2_2((~ or_tmp_37), or_tmp_23, or_191_nl);
  assign mux_33_nl = MUX_s_1_2_2(mux_32_nl, mux_29_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign weight_mem_banks_load_store_for_else_and_ssc = PECoreRun_wen & (~ mux_33_nl)
      & and_dcpl_54;
  assign nor_319_nl = ~(rva_in_reg_rw_sva_st_4 | PECore_DecodeAxiRead_switch_lp_nor_tmp_4
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 | rva_in_reg_rw_sva_4 | (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3)
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1
      | rva_in_reg_rw_sva_st_1_4);
  assign mux_64_nl = MUX_s_1_2_2(nor_319_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign weight_mem_banks_load_store_for_else_and_3_ssc = PECoreRun_wen & mux_64_nl
      & and_dcpl_54;
  assign nor_368_nl = ~((~((~(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign nor_369_nl = ~((~((~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_71_nl = MUX_s_1_2_2(nor_368_nl, nor_369_nl, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_271_nl = weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | mux_71_nl;
  assign mux_68_nl = MUX_s_1_2_2((~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])),
      (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign or_263_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]!=2'b00);
  assign mux_69_nl = MUX_s_1_2_2(mux_68_nl, or_263_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_70_nl = MUX_s_1_2_2(or_tmp_36, mux_69_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_72_nl = MUX_s_1_2_2(or_271_nl, mux_70_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_load_store_for_else_and_77_ssc = PECoreRun_wen & (~ mux_72_nl)
      & while_stage_0_6;
  assign weight_port_read_out_data_and_248_enex5 = weight_port_read_out_data_and_209_ssc
      & reg_weight_port_read_out_data_0_1_sva_dfm_1_enexo;
  assign weight_port_read_out_data_and_249_enex5 = weight_port_read_out_data_and_209_ssc
      & reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo;
  assign weight_port_read_out_data_and_250_enex5 = weight_port_read_out_data_and_209_ssc
      & reg_weight_port_read_out_data_0_2_sva_dfm_1_1_enexo;
  assign weight_port_read_out_data_and_251_enex5 = weight_port_read_out_data_and_209_ssc
      & reg_weight_port_read_out_data_0_3_sva_dfm_1_1_enexo;
  assign and_1042_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 & (~ or_dcpl_329);
  assign mux1h_9_nl = MUX1HOT_v_4_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7_4,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[7:4]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[7:4]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[7:4]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[7:4]),
      weight_port_read_out_data_0_0_sva_dfm_2_7_4, {and_1042_ssc , and_1023_cse ,
      and_1024_cse , and_1025_cse , and_1026_cse , and_1027_cse , nor_508_cse});
  assign not_2369_nl = ~ or_dcpl_329;
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w1_7_4 = MUX_v_4_2_2(4'b0000, mux1h_9_nl,
      not_2369_nl);
  assign mux1h_16_nl = MUX1HOT_v_4_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_3_0,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[3:0]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[3:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[3:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[3:0]),
      weight_port_read_out_data_0_0_sva_dfm_2_3_0, {and_1042_ssc , and_1023_cse ,
      and_1024_cse , and_1025_cse , and_1026_cse , and_1027_cse , nor_508_cse});
  assign not_2289_nl = ~ or_dcpl_329;
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w1_3_0 = MUX_v_4_2_2(4'b0000, mux1h_16_nl,
      not_2289_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_264_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_111_nl
      = MUX_v_2_2_2(2'b00, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[127:126]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_264_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_265_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_127_nl
      = MUX_v_2_2_2(2'b00, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:126]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_265_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000
      = MUX_v_2_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7_6,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1[7:6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1[7:6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1[7:6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1[7:6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1[7:6]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_111_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_127_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_145_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_128_nl
      = MUX_v_6_2_2(6'b000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[125:120]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_145_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_160_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_129_nl
      = MUX_v_6_2_2(6'b000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[125:120]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_160_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000001
      = MUX_v_6_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_5_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1[5:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_128_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_129_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_110_nl
      = (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[119]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]));
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_126_nl
      = (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[119]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000
      = MUX_s_1_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_110_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_126_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_130_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[118:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_267_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_131_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[118:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_267_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001
      = MUX_v_7_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_130_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_131_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_109_nl
      = (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[111]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]));
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_125_nl
      = (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[111]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000
      = MUX_s_1_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_109_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_125_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_132_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[110:104]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_269_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_133_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[110:104]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_269_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001
      = MUX_v_7_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_132_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_133_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign act_port_reg_data_act_port_reg_data_nor_cse = ~(PECore_RunMac_PECore_RunMac_if_and_svs_9
      | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_9));
  assign act_port_reg_data_and_16_cse = act_port_reg_data_act_port_reg_data_nor_cse
      & fsm_output;
  assign weight_port_read_out_data_and_252_enex5 = weight_port_read_out_data_and_122_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_3_enexo;
  assign weight_port_read_out_data_and_253_enex5 = weight_port_read_out_data_and_122_cse
      & reg_weight_port_read_out_data_0_2_sva_dfm_3_1_enexo;
  assign weight_port_read_out_data_and_254_enex5 = weight_port_read_out_data_and_122_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_3_1_enexo;
  assign or_33_nl = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | rva_in_reg_rw_sva_st_1_5;
  assign mux_14_nl = MUX_s_1_2_2(not_tmp_33, or_tmp_15, or_33_nl);
  assign weight_port_read_out_data_and_129_ssc = PECoreRun_wen & (~ mux_14_nl) &
      while_stage_0_7;
  assign weight_mem_run_3_for_5_and_157_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_158_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_160_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_162_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_163_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_port_read_out_data_and_130_ssc = PECoreRun_wen & ((~ mux_15_itm)
      | (~ while_stage_0_6) | PECore_RunMac_PECore_RunMac_if_and_svs_st_5) & and_dcpl_40;
  assign weight_mem_run_3_for_5_and_165_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_166_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_168_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_170_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_171_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign and_568_ssc = or_dcpl_249 & while_and_1243_cse;
  assign and_569_ssc = or_dcpl_249 & while_while_nor_259_cse;
  assign and_570_ssc = or_dcpl_249 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign nor_616_nl = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_2 | (~ mux_tmp_519));
  assign mux_552_nl = MUX_s_1_2_2(mux_tmp_519, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_553_nl = MUX_s_1_2_2(nor_616_nl, mux_552_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_554_nl = MUX_s_1_2_2(mux_tmp_519, mux_553_nl, while_stage_0_6);
  assign and_1551_cse = mux_554_nl & PECoreRun_wen;
  assign weight_port_read_out_data_and_255_enex5 = weight_port_read_out_data_and_138_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_2_enexo;
  assign weight_port_read_out_data_and_256_enex5 = weight_port_read_out_data_and_138_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo;
  assign or_1179_nl = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse
      | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse | weight_mem_run_3_for_5_and_150_itm_2
      | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse | weight_mem_run_3_for_5_and_148_itm_2
      | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse
      | weight_mem_run_3_for_5_and_cse;
  assign or_1176_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2;
  assign or_1175_nl = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2;
  assign mux_562_nl = MUX_s_1_2_2(or_1176_nl, or_1175_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign or_1174_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2;
  assign mux_563_nl = MUX_s_1_2_2(mux_562_nl, or_1174_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_1177_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1 | (crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & mux_563_nl);
  assign mux_564_nl = MUX_s_1_2_2(or_1179_nl, or_1177_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_1557_cse = mux_564_nl & weight_mem_run_3_for_aelse_and_cse;
  assign weight_port_read_out_data_and_209_ssc = PECoreRun_wen & and_dcpl_352 & while_stage_0_8
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
  assign weight_port_read_out_data_and_257_enex5 = weight_port_read_out_data_and_209_ssc
      & reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo;
  assign weight_port_read_out_data_and_258_enex5 = weight_port_read_out_data_and_209_ssc
      & reg_weight_port_read_out_data_0_0_sva_dfm_1_1_1_enexo;
  assign rva_out_reg_data_and_187_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_127_120_sva_dfm_4_1_1_enexo;
  assign rva_out_reg_data_and_188_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_119_112_sva_dfm_4_1_1_enexo;
  assign rva_out_reg_data_and_189_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_111_104_sva_dfm_4_1_1_enexo;
  assign mux_76_nl = MUX_s_1_2_2(not_tmp_33, or_tmp_15, rva_in_reg_rw_sva_st_1_5);
  assign rva_out_reg_data_and_78_ssc = PECoreRun_wen & (~ mux_76_nl) & while_stage_0_7;
  assign weight_port_read_out_data_0_1_sva_mx0_7_4 = MUX1HOT_v_4_3_2(weight_port_read_out_data_0_1_sva_dfm_1_7_4,
      weight_port_read_out_data_0_1_sva_dfm_1_1_7_4, weight_port_read_out_data_0_1_sva_7_4,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_1_sva_mx0_3_0 = MUX1HOT_v_4_3_2(weight_port_read_out_data_0_1_sva_dfm_1_3_0,
      weight_port_read_out_data_0_1_sva_dfm_1_1_3_0, weight_port_read_out_data_0_1_sva_3_0,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_7_4 = MUX1HOT_v_4_9_2(weight_port_read_out_data_0_0_sva_dfm_2_7_4,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:4]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:4]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:4]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:4]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:4]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:4]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:4]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[7:4]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse
      , weight_mem_run_3_for_5_and_148_itm_2 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse
      , weight_mem_run_3_for_5_and_150_itm_2 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_3_0 = MUX1HOT_v_4_9_2(weight_port_read_out_data_0_0_sva_dfm_2_3_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[3:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[3:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[3:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[3:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[3:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[3:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[3:0]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[3:0]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse
      , weight_mem_run_3_for_5_and_148_itm_2 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse
      , weight_mem_run_3_for_5_and_150_itm_2 , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse});
  assign weight_port_read_out_data_0_3_sva_mx0_7 = MUX1HOT_s_1_3_2(weight_port_read_out_data_0_3_sva_dfm_1_7,
      weight_port_read_out_data_0_3_sva_dfm_1_1_7, weight_port_read_out_data_0_3_sva_7,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_3_sva_mx0_6_0 = MUX1HOT_v_7_3_2(weight_port_read_out_data_0_3_sva_dfm_1_6_0,
      weight_port_read_out_data_0_3_sva_dfm_1_1_6_0, weight_port_read_out_data_0_3_sva_6_0,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_2_sva_mx0_7 = MUX1HOT_s_1_3_2(weight_port_read_out_data_0_2_sva_dfm_1_7,
      weight_port_read_out_data_0_2_sva_dfm_1_1_7, weight_port_read_out_data_0_2_sva_7,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_2_sva_mx0_6_0 = MUX1HOT_v_7_3_2(weight_port_read_out_data_0_2_sva_dfm_1_6_0,
      weight_port_read_out_data_0_2_sva_dfm_1_1_6_0, weight_port_read_out_data_0_2_sva_6_0,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign rva_out_reg_data_127_120_sva_dfm_4_mx0w0_7_6 = MUX1HOT_v_2_3_2(rva_out_reg_data_127_120_sva_dfm_7_7_6,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:126]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_35_nl = MUX_v_6_2_2(6'b000000, rva_out_reg_data_127_120_sva_dfm_6_5_0,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_127_120_sva_dfm_4_mx0w0_5_0 = MUX1HOT_v_6_3_2(while_if_while_if_and_35_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[125:120]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000001,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_119_112_sva_dfm_4_mx0w0_7 = MUX1HOT_s_1_3_2(rva_out_reg_data_119_112_sva_dfm_7_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[119]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_34_nl = MUX_v_7_2_2(7'b0000000, rva_out_reg_data_119_112_sva_dfm_6_6_0,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_119_112_sva_dfm_4_mx0w0_6_0 = MUX1HOT_v_7_3_2(while_if_while_if_and_34_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[118:112]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_111_104_sva_dfm_4_mx0w0_7 = MUX1HOT_s_1_3_2(rva_out_reg_data_111_104_sva_dfm_7_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[111]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_33_nl = MUX_v_7_2_2(7'b0000000, rva_out_reg_data_111_104_sva_dfm_6_6_0,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_111_104_sva_dfm_4_mx0w0_6_0 = MUX1HOT_v_7_3_2(while_if_while_if_and_33_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[110:104]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_and_190_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_127_120_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_191_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_119_112_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_192_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_111_104_sva_dfm_4_3_1_enexo;
  assign weight_mem_run_3_for_5_and_187_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign and_1579_nl = or_931_cse & mux_tmp_548;
  assign and_1578_nl = or_928_cse & mux_tmp_548;
  assign mux_581_nl = MUX_s_1_2_2(and_1579_nl, and_1578_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_1580_cse = mux_581_nl & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & PECoreRun_wen;
  assign and_1050_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 & (~ or_dcpl);
  assign and_1052_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      & (~ or_dcpl);
  assign and_1053_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      & (~ or_dcpl);
  assign mux1h_10_nl = MUX1HOT_v_4_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1[7:4]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[39:36]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[39:36]),
      weight_port_read_out_data_0_4_sva_mx0_7_4, {and_1050_ssc , and_1007_cse , and_1052_ssc
      , and_1053_ssc , and_1010_cse , and_1011_cse , nor_506_cse});
  assign not_2374_nl = ~ or_dcpl;
  assign weight_port_read_out_data_0_4_sva_dfm_mx0w2_7_4 = MUX_v_4_2_2(4'b0000, mux1h_10_nl,
      not_2374_nl);
  assign mux1h_17_nl = MUX1HOT_v_4_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1[3:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[35:32]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[35:32]),
      weight_port_read_out_data_0_4_sva_mx0_3_0, {and_1050_ssc , and_1007_cse , and_1052_ssc
      , and_1053_ssc , and_1010_cse , and_1011_cse , nor_506_cse});
  assign not_2291_nl = ~ or_dcpl;
  assign weight_port_read_out_data_0_4_sva_dfm_mx0w2_3_0 = MUX_v_4_2_2(4'b0000, mux1h_17_nl,
      not_2291_nl);
  assign weight_port_read_out_data_0_4_sva_mx0_7_4 = MUX1HOT_v_4_3_2(weight_port_read_out_data_0_1_sva_dfm_1_1_7_4,
      weight_port_read_out_data_0_4_sva_dfm_1_1_7_4, weight_port_read_out_data_0_4_sva_7_4,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_4_sva_mx0_3_0 = MUX1HOT_v_4_3_2(weight_port_read_out_data_0_1_sva_dfm_1_1_3_0,
      weight_port_read_out_data_0_4_sva_dfm_1_1_3_0, weight_port_read_out_data_0_4_sva_3_0,
      {and_dcpl_262 , and_dcpl_33 , (~ while_stage_0_8)});
  assign while_if_while_if_and_29_nl = MUX_v_4_2_2(4'b0000, rva_out_reg_data_87_80_sva_dfm_6_7_4,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_87_80_sva_dfm_4_mx0w0_7_4 = MUX1HOT_v_4_3_2(while_if_while_if_and_29_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:84]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_36_nl = MUX_v_4_2_2(4'b0000, rva_out_reg_data_87_80_sva_dfm_6_3_0,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_87_80_sva_dfm_4_mx0w0_3_0 = MUX1HOT_v_4_3_2(while_if_while_if_and_36_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[83:80]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000001,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_271_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_106_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[87:84]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_271_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_272_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_122_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[87:84]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_272_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000000
      = MUX_v_4_8_2(weight_port_read_out_data_0_1_sva_dfm_1_1_7_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_106_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_122_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_150_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_135_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[83:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_150_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_165_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_136_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[83:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_165_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000001
      = MUX_v_4_8_2(weight_port_read_out_data_0_1_sva_dfm_1_1_3_0, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_135_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_136_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign rva_out_reg_data_111_104_sva_dfm_7_7 = rva_out_reg_data_111_104_sva_dfm_6_7
      & rva_in_reg_rw_sva_5;
  assign rva_out_reg_data_119_112_sva_dfm_7_7 = rva_out_reg_data_119_112_sva_dfm_6_7
      & rva_in_reg_rw_sva_5;
  assign rva_out_reg_data_127_120_sva_dfm_7_7_6 = MUX_v_2_2_2(2'b00, rva_out_reg_data_127_120_sva_dfm_6_7_6,
      rva_in_reg_rw_sva_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl
      = (SC_SRAM_CONFIG[7:4]) & (signext_4_1(~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8))
      & ({{3{PECore_DecodeAxiRead_switch_lp_nor_9_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1});
  assign PECore_PushAxiRsp_if_mux1h_10_6_3 = MUX1HOT_v_4_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl,
      rva_out_reg_data_7_1_sva_dfm_6_rsp_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4[6:3]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl
      = (SC_SRAM_CONFIG[3:1]) & (signext_3_1(~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8))
      & ({{2{PECore_DecodeAxiRead_switch_lp_nor_9_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1});
  assign PECore_PushAxiRsp_if_mux1h_10_2_0 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl,
      rva_out_reg_data_7_1_sva_dfm_6_rsp_1, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4[2:0]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_20_nl = MUX_v_4_2_2((SC_SRAM_CONFIG[15:12]),
      (rva_out_reg_data_15_9_sva_dfm_9[6:3]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl
      = MUX_v_4_2_2(4'b0000, PECore_DecodeAxiRead_switch_lp_mux_20_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_12_6_3 = MUX1HOT_v_4_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl,
      rva_out_reg_data_15_9_sva_dfm_6_6_3, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4[6:3]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_6_3,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_27_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[11:9]),
      (rva_out_reg_data_15_9_sva_dfm_9[2:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl
      = MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_27_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_12_2_0 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl,
      rva_out_reg_data_15_9_sva_dfm_6_2_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4[2:0]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_2_0,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_21_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[23]),
      (rva_out_reg_data_23_17_sva_dfm_7[6]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl
      = PECore_DecodeAxiRead_switch_lp_mux_21_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_14_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl,
      rva_out_reg_data_23_17_sva_dfm_6_6, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4[6]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_6, {PECore_PushAxiRsp_if_asn_79
      , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_28_nl = MUX_v_6_2_2((SC_SRAM_CONFIG[22:17]),
      (rva_out_reg_data_23_17_sva_dfm_7[5:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl
      = MUX_v_6_2_2(6'b000000, PECore_DecodeAxiRead_switch_lp_mux_28_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_14_5_0 = MUX1HOT_v_6_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl,
      rva_out_reg_data_23_17_sva_dfm_6_5_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4[5:0]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_5_0,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign rva_out_reg_data_and_193_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_194_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_195_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_196_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_197_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_198_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_1_1_enexo;
  assign rva_out_reg_data_and_199_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_200_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_1_1_enexo;
  assign or_tmp_484 = PECore_UpdateFSM_switch_lp_equal_tmp_2_9 | act_port_reg_data_act_port_reg_data_nor_cse;
  assign not_tmp_488 = ~(while_stage_0_10 | (~ or_tmp_484));
  assign or_929_nl = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2_cse
      | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_2 | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse
      | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse;
  assign mux_tmp_427 = MUX_s_1_2_2(or_dcpl_243, or_929_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign or_933_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
      | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2 | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse
      | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse;
  assign mux_tmp_429 = MUX_s_1_2_2(or_dcpl_243, or_933_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign and_dcpl_949 = while_stage_0_3 & fsm_output;
  assign and_dcpl_958 = fsm_output & while_stage_0_7;
  assign or_dcpl_390 = weight_mem_run_3_for_5_and_31_itm_2 | weight_mem_run_3_for_5_and_142_itm_1;
  assign or_dcpl_394 = weight_mem_run_3_for_5_and_30_itm_2 | weight_mem_run_3_for_5_and_28_itm_2;
  assign or_dcpl_395 = weight_mem_run_3_for_5_and_136_itm_1 | weight_mem_run_3_for_5_and_135_itm_1;
  assign or_dcpl_403 = weight_mem_run_3_for_5_and_135_itm_1 | weight_mem_run_3_for_5_and_30_itm_2;
  assign or_dcpl_407 = weight_mem_run_3_for_5_and_142_itm_1 | weight_mem_run_3_for_5_and_28_itm_2;
  assign or_dcpl_408 = weight_mem_run_3_for_5_and_136_itm_1 | weight_mem_run_3_for_5_and_31_itm_2;
  assign or_tmp_541 = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  assign mux_492_nl = MUX_s_1_2_2((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]),
      (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])), reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign mux_493_nl = MUX_s_1_2_2(mux_492_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_1054_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | mux_493_nl;
  assign mux_494_cse = MUX_s_1_2_2(nand_76_cse, or_1054_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_tmp_17 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7 & (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 | mux_494_cse);
  assign and_tmp_18 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7 & (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 | mux_494_cse);
  assign or_1122_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1;
  assign or_1121_nl = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1;
  assign mux_520_nl = MUX_s_1_2_2(or_1122_nl, or_1121_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign or_1120_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1;
  assign mux_521_nl = MUX_s_1_2_2(mux_520_nl, or_1120_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_tmp_583 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | mux_521_nl;
  assign or_tmp_584 = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | rva_in_reg_rw_sva_st_1_5 | (~ or_tmp_583);
  assign or_1125_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      | (~ while_stage_0_8) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1;
  assign mux_522_cse = MUX_s_1_2_2(or_1125_nl, or_tmp_583, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign or_1146_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1;
  assign or_1145_nl = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1;
  assign mux_538_nl = MUX_s_1_2_2(or_1146_nl, or_1145_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign or_1144_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1;
  assign mux_539_nl = MUX_s_1_2_2(mux_538_nl, or_1144_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_tmp_607 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | mux_539_nl;
  assign or_tmp_608 = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | rva_in_reg_rw_sva_st_1_5 | (~ or_tmp_607);
  assign or_1149_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      | (~ while_stage_0_8) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1;
  assign mux_540_itm = MUX_s_1_2_2(or_1149_nl, or_tmp_607, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign or_1151_nl = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2;
  assign mux_tmp_512 = MUX_s_1_2_2(or_dcpl_243, or_1151_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign or_1155_nl = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2;
  assign mux_tmp_514 = MUX_s_1_2_2(or_dcpl_243, or_1155_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign and_1626_nl = ((~ while_stage_0_8) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
      | weight_mem_run_3_for_land_1_lpi_1_dfm_3) & while_stage_0_7;
  assign and_1627_nl = ((~ while_stage_0_8) | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1)
      & while_stage_0_7;
  assign and_1628_nl = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1)
      & while_stage_0_7;
  assign and_1629_nl = ((~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1)
      & while_stage_0_7;
  assign mux_548_nl = MUX_s_1_2_2(and_1628_nl, and_1629_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign and_1630_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1)
      & while_stage_0_7;
  assign mux_549_nl = MUX_s_1_2_2(mux_548_nl, and_1630_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign mux_550_nl = MUX_s_1_2_2(and_1627_nl, mux_549_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign mux_tmp_519 = MUX_s_1_2_2(and_1626_nl, mux_550_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_1204_nl = reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2_cse
      | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2;
  assign mux_tmp_548 = MUX_s_1_2_2(or_dcpl_243, or_1204_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign data_in_tmp_operator_2_for_and_15_tmp = PECoreRun_wen & and_dcpl_40 & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign data_in_tmp_operator_2_for_and_31_tmp = PECoreRun_wen & and_dcpl_40 & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign pe_manager_base_input_and_tmp = PECoreRun_wen & ((nand_91_cse & while_stage_0_3)
      | and_cse);
  assign rva_in_reg_data_and_tmp = PECoreRun_wen & and_dcpl_314 & (and_315_cse |
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign input_mem_banks_read_1_read_data_and_4_tmp = PECoreRun_wen & (while_and_4_cse
      | ((~ reg_rva_in_reg_rw_sva_st_1_1_cse) & ProductSum_for_asn_56_itm_1 & and_dcpl_205));
  assign or_1051_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~((~ while_stage_0_3)
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 | (~(reg_rva_in_reg_rw_sva_st_1_1_cse
      & ((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:0]!=16'b0000000000000001)) &
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt))));
  assign mux_491_nl = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, or_1051_nl,
      nor_524_cse);
  assign and_1434_tmp = (~ mux_491_nl) & and_cse & PECoreRun_wen;
  assign mux_542_nl = MUX_s_1_2_2((~ mux_540_itm), or_tmp_608, and_1607_cse);
  assign mux_541_nl = MUX_s_1_2_2((~ mux_540_itm), or_tmp_608, and_1608_cse);
  assign mux_543_nl = MUX_s_1_2_2(mux_542_nl, mux_541_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_1538_tmp = (~ mux_543_nl) & and_dcpl_47 & PECoreRun_wen;
  assign accum_vector_data_and_55_cse = while_stage_0_10 & fsm_output;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_cgo_ir_cse <=
          1'b0;
      reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_cgo_ir_cse <=
          1'b0;
      reg_PECore_RunScale_if_for_4_mul_1_cmp_cgo_ir_7_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_act_port_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      weight_port_read_out_data_7_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_9_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_11_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_10_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_13_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_12_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_15_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_14_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_15_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_14_sva_dfm_1 <= 8'b00000000;
      pe_config_manager_counter_sva_dfm_3_1 <= 4'b0000;
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= 1'b0;
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= 1'b0;
      while_stage_0_3 <= 1'b0;
      while_stage_0_4 <= 1'b0;
      while_stage_0_5 <= 1'b0;
      while_stage_0_6 <= 1'b0;
      while_stage_0_7 <= 1'b0;
      while_stage_0_8 <= 1'b0;
      while_stage_0_9 <= 1'b0;
      while_stage_0_10 <= 1'b0;
      while_stage_0_11 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1
          <= 1'b0;
      input_read_addrs_sva_1_1 <= 8'b00000000;
      ProductSum_for_asn_56_itm_1 <= 1'b0;
      ProductSum_for_asn_82_itm_1 <= 1'b0;
      ProductSum_for_asn_69_itm_1 <= 1'b0;
      ProductSum_for_asn_95_itm_1 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1 <= 1'b0;
      PECore_RunMac_PECore_RunMac_if_and_svs_1 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1 <= 1'b0;
      weight_port_read_out_data_0_3_sva_7 <= 1'b0;
      weight_port_read_out_data_0_2_sva_7 <= 1'b0;
    end
    else if ( PECoreRun_wen ) begin
      reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_cgo_ir_cse <=
          and_511_rmff;
      reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_cgo_ir_cse <=
          and_514_rmff;
      reg_PECore_RunScale_if_for_4_mul_1_cmp_cgo_ir_7_cse <= and_516_rmff;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= and_520_rmff;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= and_523_rmff;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= and_527_rmff;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= and_531_rmff;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= and_534_rmff;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= and_537_rmff;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= and_540_rmff;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= and_543_rmff;
      reg_rva_out_Push_mioi_iswt0_cse <= and_545_cse;
      reg_start_PopNB_mioi_iswt0_cse <= and_547_rmff;
      reg_act_port_Push_mioi_iswt0_cse <= and_549_cse;
      reg_rva_in_PopNB_mioi_iswt0_cse <= fsm_output;
      weight_port_read_out_data_7_0_sva_dfm_1 <= weight_port_read_out_data_7_0_sva_dfm_1_2;
      weight_port_read_out_data_7_3_sva_dfm_1 <= weight_port_read_out_data_7_3_sva_dfm_1_2;
      weight_port_read_out_data_7_2_sva_dfm_1 <= weight_port_read_out_data_7_2_sva_dfm_1_2;
      weight_port_read_out_data_7_5_sva_dfm_1 <= weight_port_read_out_data_7_5_sva_dfm_1_2;
      weight_port_read_out_data_7_4_sva_dfm_1 <= weight_port_read_out_data_7_4_sva_dfm_1_2;
      weight_port_read_out_data_7_7_sva_dfm_1 <= weight_port_read_out_data_7_7_sva_dfm_1_2;
      weight_port_read_out_data_7_6_sva_dfm_1 <= weight_port_read_out_data_7_6_sva_dfm_1_2;
      weight_port_read_out_data_7_9_sva_dfm_1 <= weight_port_read_out_data_7_9_sva_dfm_1_2;
      weight_port_read_out_data_7_8_sva_dfm_1 <= weight_port_read_out_data_7_8_sva_dfm_1_2;
      weight_port_read_out_data_7_11_sva_dfm_1 <= weight_port_read_out_data_7_11_sva_dfm_1_2;
      weight_port_read_out_data_7_10_sva_dfm_1 <= weight_port_read_out_data_7_10_sva_dfm_1_2;
      weight_port_read_out_data_7_13_sva_dfm_1 <= weight_port_read_out_data_7_13_sva_dfm_1_2;
      weight_port_read_out_data_7_12_sva_dfm_1 <= weight_port_read_out_data_7_12_sva_dfm_1_2;
      weight_port_read_out_data_7_15_sva_dfm_1 <= weight_port_read_out_data_7_15_sva_dfm_1_2;
      weight_port_read_out_data_7_14_sva_dfm_1 <= weight_port_read_out_data_7_14_sva_dfm_1_2;
      weight_port_read_out_data_5_15_sva_dfm_1 <= weight_port_read_out_data_5_15_sva_dfm_1_2;
      weight_port_read_out_data_5_14_sva_dfm_1 <= weight_port_read_out_data_5_14_sva_dfm_1_2;
      pe_config_manager_counter_sva_dfm_3_1 <= MUX_v_4_2_2(4'b0000, operator_4_false_acc_nl,
          pe_config_UpdateManagerCounter_if_not_7_nl);
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= ~((pe_config_input_counter_sva_mx1 != (operator_16_false_acc_sdt_sva_1[7:0]))
          | (operator_16_false_acc_sdt_sva_1[8]));
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
      while_stage_0_3 <= reg_rva_in_PopNB_mioi_iswt0_cse;
      while_stage_0_4 <= while_stage_0_3;
      while_stage_0_5 <= while_stage_0_4;
      while_stage_0_6 <= while_stage_0_5;
      while_stage_0_7 <= while_stage_0_6;
      while_stage_0_8 <= while_stage_0_7;
      while_stage_0_9 <= while_stage_0_8;
      while_stage_0_10 <= while_stage_0_9;
      while_stage_0_11 <= while_stage_0_10;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1 <= ~ (pe_manager_base_weight_sva_mx2[1]);
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 <= pe_manager_base_weight_sva_mx3_0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1 <= pe_manager_base_weight_sva_mx2[1];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[2];
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= (pe_manager_base_weight_sva_mx1_3_0[2])
          & pe_manager_base_weight_sva_mx3_0 & (~ (pe_manager_base_weight_sva_mx2[1]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1
          <= ~((pe_manager_base_weight_sva_mx1_3_0[2]) | (pe_manager_base_weight_sva_mx2[1])
          | pe_manager_base_weight_sva_mx3_0);
      input_read_addrs_sva_1_1 <= nl_input_read_addrs_sva_1_1[7:0];
      ProductSum_for_asn_56_itm_1 <= MUX1HOT_s_1_3_2(accum_vector_data_5_sva_1_load_mx0w0,
          accum_vector_data_5_sva_1_load, input_read_req_valid_lpi_1_dfm_1_mx0w2,
          {and_dcpl_658 , and_dcpl_659 , rva_in_PopNB_mioi_return_rsc_z_mxwt});
      ProductSum_for_asn_82_itm_1 <= MUX_s_1_2_2(accum_vector_data_3_sva_1_load_mx0w1,
          accum_vector_data_3_sva_1_load, or_dcpl_259);
      ProductSum_for_asn_69_itm_1 <= MUX1HOT_s_1_3_2(accum_vector_data_4_sva_1_load_mx0w0,
          accum_vector_data_4_sva_1_load, input_read_req_valid_lpi_1_dfm_1_mx0w2,
          {and_dcpl_658 , and_dcpl_659 , rva_in_PopNB_mioi_return_rsc_z_mxwt});
      ProductSum_for_asn_95_itm_1 <= MUX_s_1_2_2(accum_vector_data_2_sva_1_load_mx0w0,
          accum_vector_data_2_sva_1_load, or_dcpl_259);
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_1 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= MUX1HOT_s_1_3_2(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_mx0w0,
          accum_vector_data_0_sva_1_load_mx0w1, accum_vector_data_0_sva_1_load, {rva_in_PopNB_mioi_return_rsc_z_mxwt
          , and_dcpl_658 , and_dcpl_659});
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1 <= MUX1HOT_s_1_3_2(and_315_cse,
          accum_vector_data_1_sva_1_load_mx0w1, accum_vector_data_1_sva_1_load, {rva_in_PopNB_mioi_return_rsc_z_mxwt
          , and_dcpl_658 , and_dcpl_659});
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1 <= MUX1HOT_s_1_3_2(PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0,
          accum_vector_data_7_sva_1_load_mx0w1, accum_vector_data_7_sva_1_load, {rva_in_PopNB_mioi_return_rsc_z_mxwt
          , and_dcpl_658 , and_dcpl_659});
      PECore_RunMac_PECore_RunMac_if_and_svs_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1 <= MUX1HOT_s_1_3_2(PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0,
          accum_vector_data_6_sva_1_load_mx0w1, accum_vector_data_6_sva_1_load, {rva_in_PopNB_mioi_return_rsc_z_mxwt
          , and_dcpl_658 , and_dcpl_659});
      weight_port_read_out_data_0_3_sva_7 <= weight_port_read_out_data_0_3_sva_mx0_7;
      weight_port_read_out_data_0_2_sva_7 <= weight_port_read_out_data_0_2_sva_mx0_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_2_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_128_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= rva_out_reg_data_15_9_sva_dfm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_7 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_129_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_7 <= rva_out_reg_data_23_17_sva_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_130_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= rva_out_reg_data_30_25_sva_dfm_6_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_131_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd <= rva_out_reg_data_103_96_sva_dfm_4_3_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_132_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_103_96_sva_dfm_4_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_88_sva_dfm_4_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_133_enex5 ) begin
      rva_out_reg_data_95_88_sva_dfm_4_4 <= rva_out_reg_data_95_88_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_4_ftd <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_134_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_4_ftd <= rva_out_reg_data_87_80_sva_dfm_4_3_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_4_ftd_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_135_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_87_80_sva_dfm_4_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_72_sva_dfm_4_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_136_enex5 ) begin
      rva_out_reg_data_79_72_sva_dfm_4_4 <= rva_out_reg_data_79_72_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_4_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_137_enex5 ) begin
      rva_out_reg_data_71_64_sva_dfm_4_4 <= rva_out_reg_data_71_64_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_63_sva_dfm_4_4 <= 1'b0;
      rva_out_reg_data_47_sva_dfm_4_4 <= 1'b0;
      input_read_req_valid_lpi_1_dfm_1_9 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= 1'b0;
      rva_out_reg_data_127_120_sva_dfm_4_4_7_6 <= 2'b00;
      rva_out_reg_data_119_112_sva_dfm_4_4_7 <= 1'b0;
      rva_out_reg_data_111_104_sva_dfm_4_4_7 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_26_cse ) begin
      rva_out_reg_data_63_sva_dfm_4_4 <= PECore_RunMac_PECore_RunMac_if_and_svs_8;
      rva_out_reg_data_47_sva_dfm_4_4 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      input_read_req_valid_lpi_1_dfm_1_9 <= input_read_req_valid_lpi_1_dfm_1_8;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
      rva_out_reg_data_127_120_sva_dfm_4_4_7_6 <= reg_rva_out_reg_data_127_120_sva_dfm_4_3_ftd;
      rva_out_reg_data_119_112_sva_dfm_4_4_7 <= reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd;
      rva_out_reg_data_111_104_sva_dfm_4_4_7 <= reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_138_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_4 <= rva_out_reg_data_62_56_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_139_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= rva_out_reg_data_35_32_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_140_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_4 <= rva_out_reg_data_55_48_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_141_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_4 <= rva_out_reg_data_39_36_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_142_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_4 <= rva_out_reg_data_46_40_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1 <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1
          <= 3'b000;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_2_0 <=
          3'b000;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_6 <=
          1'b0;
      weight_port_read_out_data_0_3_sva_dfm_4_7 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_122_cse ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1 <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1[0];
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1
          <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1[3:1];
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1 <= reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1[0];
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1 <= reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_1[0];
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_2_0 <=
          reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1[3:1];
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_6 <=
          reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd;
      weight_port_read_out_data_0_3_sva_dfm_4_7 <= reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_35_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd
          <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_213_enex5 ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd
          <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_36_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_37_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_6 <= 6'b000000;
      rva_out_reg_data_0_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_8_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_16_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_31_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_24_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_0 <= 4'b0000;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_1 <= 3'b000;
      rva_out_reg_data_15_9_sva_dfm_6_6_3 <= 4'b0000;
      rva_out_reg_data_15_9_sva_dfm_6_2_0 <= 3'b000;
      rva_out_reg_data_23_17_sva_dfm_6_6 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_6_5_0 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_16;
      rva_out_reg_data_0_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_24_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
      rva_out_reg_data_8_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_25_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
      rva_out_reg_data_16_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_26_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
      rva_out_reg_data_31_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_17;
      rva_out_reg_data_24_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_15;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_0 <= PECore_PushAxiRsp_if_mux1h_10_6_3;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_1 <= PECore_PushAxiRsp_if_mux1h_10_2_0;
      rva_out_reg_data_15_9_sva_dfm_6_6_3 <= PECore_PushAxiRsp_if_mux1h_12_6_3;
      rva_out_reg_data_15_9_sva_dfm_6_2_0 <= PECore_PushAxiRsp_if_mux1h_12_2_0;
      rva_out_reg_data_23_17_sva_dfm_6_6 <= PECore_PushAxiRsp_if_mux1h_14_6;
      rva_out_reg_data_23_17_sva_dfm_6_5_0 <= PECore_PushAxiRsp_if_mux1h_14_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_38_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_9 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_cse ) begin
      rva_in_reg_rw_sva_9 <= rva_in_reg_rw_sva_8;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_9 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_6 ) begin
      rva_in_reg_rw_sva_st_1_9 <= rva_in_reg_rw_sva_st_1_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= 1'b0;
    end
    else if ( PECore_PushOutput_if_and_cse ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_27_0_sva <= 28'b0000000000000000000000000000;
      act_port_reg_data_59_32_sva <= 28'b0000000000000000000000000000;
      act_port_reg_data_91_64_sva <= 28'b0000000000000000000000000000;
      act_port_reg_data_123_96_sva <= 28'b0000000000000000000000000000;
      act_port_reg_data_155_128_sva <= 28'b0000000000000000000000000000;
      act_port_reg_data_187_160_sva <= 28'b0000000000000000000000000000;
      act_port_reg_data_219_192_sva <= 28'b0000000000000000000000000000;
      act_port_reg_data_251_224_sva <= 28'b0000000000000000000000000000;
    end
    else if ( and_1086_cse ) begin
      act_port_reg_data_27_0_sva <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (PECore_RunScale_if_for_4_mul_1_cmp_2_z[38:11]), PECore_UpdateFSM_switch_lp_not_23_nl);
      act_port_reg_data_59_32_sva <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (PECore_RunScale_if_for_4_mul_1_cmp_4_z[38:11]), PECore_UpdateFSM_switch_lp_not_24_nl);
      act_port_reg_data_91_64_sva <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (PECore_RunScale_if_for_4_mul_1_cmp_6_z[38:11]), PECore_UpdateFSM_switch_lp_not_25_nl);
      act_port_reg_data_123_96_sva <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (PECore_RunScale_if_for_4_mul_1_cmp_z[38:11]), PECore_UpdateFSM_switch_lp_not_26_nl);
      act_port_reg_data_155_128_sva <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (PECore_RunScale_if_for_4_mul_1_cmp_7_z[38:11]), PECore_UpdateFSM_switch_lp_not_27_nl);
      act_port_reg_data_187_160_sva <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (PECore_RunScale_if_for_4_mul_1_cmp_5_z[38:11]), PECore_UpdateFSM_switch_lp_not_28_nl);
      act_port_reg_data_219_192_sva <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (PECore_RunScale_if_for_4_mul_1_cmp_3_z[38:11]), PECore_UpdateFSM_switch_lp_not_29_nl);
      act_port_reg_data_251_224_sva <= MUX_v_28_2_2(28'b0000000000000000000000000000,
          (PECore_RunScale_if_for_4_mul_1_cmp_1_z[38:11]), PECore_UpdateFSM_switch_lp_not_19_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= 1'b0;
      PECore_RunMac_PECore_RunMac_if_and_svs_9 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
      PECore_RunMac_PECore_RunMac_if_and_svs_9 <= PECore_RunMac_PECore_RunMac_if_and_svs_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_sva <= 31'b0000000000000000000000000000000;
      accum_vector_data_6_sva <= 31'b0000000000000000000000000000000;
      accum_vector_data_5_sva <= 31'b0000000000000000000000000000000;
      accum_vector_data_4_sva <= 31'b0000000000000000000000000000000;
      accum_vector_data_3_sva <= 31'b0000000000000000000000000000000;
      accum_vector_data_2_sva <= 31'b0000000000000000000000000000000;
      accum_vector_data_1_sva <= 31'b0000000000000000000000000000000;
      accum_vector_data_0_sva <= 31'b0000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_cse ) begin
      accum_vector_data_7_sva <= accum_vector_data_acc_itm;
      accum_vector_data_6_sva <= accum_vector_data_acc_26_itm;
      accum_vector_data_5_sva <= accum_vector_data_acc_23_itm;
      accum_vector_data_4_sva <= accum_vector_data_acc_20_itm;
      accum_vector_data_3_sva <= accum_vector_data_acc_17_itm;
      accum_vector_data_2_sva <= accum_vector_data_acc_14_itm;
      accum_vector_data_1_sva <= accum_vector_data_acc_11_itm;
      accum_vector_data_0_sva <= accum_vector_data_acc_8_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_8 <= 1'b0;
      rva_in_reg_rw_sva_st_8 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_2_cse ) begin
      rva_in_reg_rw_sva_st_1_8 <= rva_in_reg_rw_sva_st_1_7;
      rva_in_reg_rw_sva_st_8 <= rva_in_reg_rw_sva_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_sva_8 <= 31'b0000000000000000000000000000000;
      accum_vector_data_7_sva_7 <= 31'b0000000000000000000000000000000;
      accum_vector_data_7_sva_6 <= 31'b0000000000000000000000000000000;
      accum_vector_data_7_sva_5 <= 31'b0000000000000000000000000000000;
      accum_vector_data_7_sva_4 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1125_cse ) begin
      accum_vector_data_7_sva_8 <= accum_vector_data_7_sva_8_mx0w0;
      accum_vector_data_7_sva_7 <= accum_vector_data_7_sva_7_mx0w0;
      accum_vector_data_7_sva_6 <= accum_vector_data_7_sva_6_mx0w0;
      accum_vector_data_7_sva_5 <= accum_vector_data_7_sva_5_mx0w0;
      accum_vector_data_7_sva_4 <= accum_vector_data_7_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_6_sva_8 <= 31'b0000000000000000000000000000000;
      accum_vector_data_6_sva_7 <= 31'b0000000000000000000000000000000;
      accum_vector_data_6_sva_6 <= 31'b0000000000000000000000000000000;
      accum_vector_data_6_sva_5 <= 31'b0000000000000000000000000000000;
      accum_vector_data_6_sva_4 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1140_cse ) begin
      accum_vector_data_6_sva_8 <= accum_vector_data_6_sva_8_mx0w0;
      accum_vector_data_6_sva_7 <= accum_vector_data_6_sva_7_mx0w0;
      accum_vector_data_6_sva_6 <= accum_vector_data_6_sva_6_mx0w0;
      accum_vector_data_6_sva_5 <= accum_vector_data_6_sva_5_mx0w0;
      accum_vector_data_6_sva_4 <= accum_vector_data_6_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_5_sva_8 <= 31'b0000000000000000000000000000000;
      accum_vector_data_5_sva_7 <= 31'b0000000000000000000000000000000;
      accum_vector_data_5_sva_6 <= 31'b0000000000000000000000000000000;
      accum_vector_data_5_sva_5 <= 31'b0000000000000000000000000000000;
      accum_vector_data_5_sva_4 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1155_cse ) begin
      accum_vector_data_5_sva_8 <= accum_vector_data_5_sva_8_mx0w0;
      accum_vector_data_5_sva_7 <= accum_vector_data_5_sva_7_mx0w0;
      accum_vector_data_5_sva_6 <= accum_vector_data_5_sva_6_mx0w0;
      accum_vector_data_5_sva_5 <= accum_vector_data_5_sva_5_mx0w0;
      accum_vector_data_5_sva_4 <= accum_vector_data_5_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_4_sva_9 <= 31'b0000000000000000000000000000000;
      accum_vector_data_4_sva_8 <= 31'b0000000000000000000000000000000;
      accum_vector_data_4_sva_7 <= 31'b0000000000000000000000000000000;
      accum_vector_data_4_sva_6 <= 31'b0000000000000000000000000000000;
      accum_vector_data_4_sva_5 <= 31'b0000000000000000000000000000000;
      accum_vector_data_4_sva_4 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1170_cse ) begin
      accum_vector_data_4_sva_9 <= accum_vector_data_4_sva_9_mx0w0;
      accum_vector_data_4_sva_8 <= accum_vector_data_4_sva_8_mx0w0;
      accum_vector_data_4_sva_7 <= accum_vector_data_4_sva_7_mx0w0;
      accum_vector_data_4_sva_6 <= accum_vector_data_4_sva_6_mx0w0;
      accum_vector_data_4_sva_5 <= accum_vector_data_4_sva_5_mx0w0;
      accum_vector_data_4_sva_4 <= accum_vector_data_4_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_3_sva_8 <= 31'b0000000000000000000000000000000;
      accum_vector_data_3_sva_7 <= 31'b0000000000000000000000000000000;
      accum_vector_data_3_sva_6 <= 31'b0000000000000000000000000000000;
      accum_vector_data_3_sva_5 <= 31'b0000000000000000000000000000000;
      accum_vector_data_3_sva_4 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1188_cse ) begin
      accum_vector_data_3_sva_8 <= accum_vector_data_3_sva_8_mx0w0;
      accum_vector_data_3_sva_7 <= accum_vector_data_3_sva_7_mx0w0;
      accum_vector_data_3_sva_6 <= accum_vector_data_3_sva_6_mx0w0;
      accum_vector_data_3_sva_5 <= accum_vector_data_3_sva_5_mx0w0;
      accum_vector_data_3_sva_4 <= accum_vector_data_3_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_2_sva_9 <= 31'b0000000000000000000000000000000;
      accum_vector_data_2_sva_8 <= 31'b0000000000000000000000000000000;
      accum_vector_data_2_sva_7 <= 31'b0000000000000000000000000000000;
      accum_vector_data_2_sva_6 <= 31'b0000000000000000000000000000000;
      accum_vector_data_2_sva_5 <= 31'b0000000000000000000000000000000;
      accum_vector_data_2_sva_4 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1203_cse ) begin
      accum_vector_data_2_sva_9 <= accum_vector_data_2_sva_9_mx0w0;
      accum_vector_data_2_sva_8 <= accum_vector_data_2_sva_8_mx0w0;
      accum_vector_data_2_sva_7 <= accum_vector_data_2_sva_7_mx0w0;
      accum_vector_data_2_sva_6 <= accum_vector_data_2_sva_6_mx0w0;
      accum_vector_data_2_sva_5 <= accum_vector_data_2_sva_5_mx0w0;
      accum_vector_data_2_sva_4 <= accum_vector_data_2_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_1_sva_8 <= 31'b0000000000000000000000000000000;
      accum_vector_data_1_sva_7 <= 31'b0000000000000000000000000000000;
      accum_vector_data_1_sva_6 <= 31'b0000000000000000000000000000000;
      accum_vector_data_1_sva_5 <= 31'b0000000000000000000000000000000;
      accum_vector_data_1_sva_4 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1221_cse ) begin
      accum_vector_data_1_sva_8 <= accum_vector_data_1_sva_8_mx0w0;
      accum_vector_data_1_sva_7 <= accum_vector_data_1_sva_7_mx0w0;
      accum_vector_data_1_sva_6 <= accum_vector_data_1_sva_6_mx0w0;
      accum_vector_data_1_sva_5 <= accum_vector_data_1_sva_5_mx0w0;
      accum_vector_data_1_sva_4 <= accum_vector_data_1_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_0_sva_8 <= 31'b0000000000000000000000000000000;
      accum_vector_data_0_sva_7 <= 31'b0000000000000000000000000000000;
      accum_vector_data_0_sva_6 <= 31'b0000000000000000000000000000000;
      accum_vector_data_0_sva_5 <= 31'b0000000000000000000000000000000;
      accum_vector_data_0_sva_4 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1236_cse ) begin
      accum_vector_data_0_sva_8 <= accum_vector_data_0_sva_8_mx0w0;
      accum_vector_data_0_sva_7 <= accum_vector_data_0_sva_7_mx0w0;
      accum_vector_data_0_sva_6 <= accum_vector_data_0_sva_6_mx0w0;
      accum_vector_data_0_sva_5 <= accum_vector_data_0_sva_5_mx0w0;
      accum_vector_data_0_sva_4 <= accum_vector_data_0_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_29 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_7)
        ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_operator_1_for_asn_115_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_100_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_85_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_73_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_55_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_43_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_25_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_10_itm_7 <= 1'b0;
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= 1'b0;
    end
    else if ( accum_vector_operator_1_for_and_cse ) begin
      accum_vector_operator_1_for_asn_115_itm_7 <= accum_vector_operator_1_for_asn_118_itm_6;
      accum_vector_operator_1_for_asn_100_itm_7 <= accum_vector_operator_1_for_asn_103_itm_6;
      accum_vector_operator_1_for_asn_85_itm_7 <= accum_vector_operator_1_for_asn_88_itm_6;
      accum_vector_operator_1_for_asn_73_itm_7 <= accum_vector_operator_1_for_asn_73_itm_6;
      accum_vector_operator_1_for_asn_55_itm_7 <= accum_vector_operator_1_for_asn_58_itm_6;
      accum_vector_operator_1_for_asn_43_itm_7 <= accum_vector_operator_1_for_asn_43_itm_6;
      accum_vector_operator_1_for_asn_25_itm_7 <= accum_vector_operator_1_for_asn_28_itm_6;
      accum_vector_operator_1_for_asn_10_itm_7 <= accum_vector_operator_1_for_asn_13_itm_6;
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_sva_9 <= 31'b0000000000000000000000000000000;
    end
    else if ( while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
        & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_118_itm_6)
        ) begin
      accum_vector_data_7_sva_9 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ProductSum_for_acc_20_cmp_z, accum_vector_operator_1_for_not_39_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_6_sva_9 <= 31'b0000000000000000000000000000000;
    end
    else if ( while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
        & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_103_itm_6)
        ) begin
      accum_vector_data_6_sva_9 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_z, accum_vector_operator_1_for_not_38_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_5_sva_9 <= 31'b0000000000000000000000000000000;
    end
    else if ( while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
        & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_88_itm_6)
        ) begin
      accum_vector_data_5_sva_9 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_z, accum_vector_operator_1_for_not_37_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_3_sva_9 <= 31'b0000000000000000000000000000000;
    end
    else if ( while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
        & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_58_itm_6)
        ) begin
      accum_vector_data_3_sva_9 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_z, accum_vector_operator_1_for_not_36_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_1_sva_9 <= 31'b0000000000000000000000000000000;
    end
    else if ( while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
        & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_28_itm_6)
        ) begin
      accum_vector_data_1_sva_9 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_z, accum_vector_operator_1_for_not_35_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_0_sva_9 <= 31'b0000000000000000000000000000000;
    end
    else if ( while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
        & PECoreRun_wen & (PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_13_itm_6)
        ) begin
      accum_vector_data_0_sva_9 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_z, accum_vector_operator_1_for_not_34_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= 1'b0;
      rva_in_reg_rw_sva_8 <= 1'b0;
    end
    else if ( while_if_and_6_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
      rva_in_reg_rw_sva_8 <= rva_in_reg_rw_sva_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
        | PECore_RunMac_PECore_RunMac_if_and_svs_st_6)) & while_stage_0_8 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= 1'b0;
      accum_vector_operator_1_for_asn_118_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_103_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_88_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_58_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_28_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_13_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_73_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_43_itm_6 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_2_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
      accum_vector_operator_1_for_asn_118_itm_6 <= accum_vector_operator_1_for_asn_118_itm_5;
      accum_vector_operator_1_for_asn_103_itm_6 <= accum_vector_operator_1_for_asn_103_itm_5;
      accum_vector_operator_1_for_asn_88_itm_6 <= accum_vector_operator_1_for_asn_88_itm_5;
      accum_vector_operator_1_for_asn_58_itm_6 <= accum_vector_operator_1_for_asn_58_itm_5;
      accum_vector_operator_1_for_asn_28_itm_6 <= accum_vector_operator_1_for_asn_28_itm_5;
      accum_vector_operator_1_for_asn_13_itm_6 <= accum_vector_operator_1_for_asn_13_itm_5;
      accum_vector_operator_1_for_asn_73_itm_6 <= accum_vector_operator_1_for_asn_73_itm_5;
      accum_vector_operator_1_for_asn_43_itm_6 <= accum_vector_operator_1_for_asn_43_itm_5;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= 1'b0;
      weight_port_read_out_data_0_7_sva <= 8'b00000000;
      weight_port_read_out_data_0_5_sva <= 8'b00000000;
      rva_in_reg_rw_sva_7 <= 1'b0;
      weight_port_read_out_data_0_1_sva_7_4 <= 4'b0000;
      weight_port_read_out_data_0_1_sva_3_0 <= 4'b0000;
      weight_port_read_out_data_0_3_sva_6_0 <= 7'b0000000;
      weight_port_read_out_data_0_2_sva_6_0 <= 7'b0000000;
      weight_port_read_out_data_0_4_sva_7_4 <= 4'b0000;
      weight_port_read_out_data_0_4_sva_3_0 <= 4'b0000;
    end
    else if ( while_if_and_7_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6;
      weight_port_read_out_data_0_7_sva <= weight_port_read_out_data_0_7_sva_mx0;
      weight_port_read_out_data_0_5_sva <= weight_port_read_out_data_0_5_sva_mx0;
      rva_in_reg_rw_sva_7 <= rva_in_reg_rw_sva_6;
      weight_port_read_out_data_0_1_sva_7_4 <= weight_port_read_out_data_0_1_sva_mx0_7_4;
      weight_port_read_out_data_0_1_sva_3_0 <= weight_port_read_out_data_0_1_sva_mx0_3_0;
      weight_port_read_out_data_0_3_sva_6_0 <= weight_port_read_out_data_0_3_sva_mx0_6_0;
      weight_port_read_out_data_0_2_sva_6_0 <= weight_port_read_out_data_0_2_sva_mx0_6_0;
      weight_port_read_out_data_0_4_sva_7_4 <= weight_port_read_out_data_0_4_sva_mx0_7_4;
      weight_port_read_out_data_0_4_sva_3_0 <= weight_port_read_out_data_0_4_sva_mx0_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_26_itm_6 <= 1'b0;
      ProductSum_for_asn_40_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_96_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_99_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_98_itm_1 <= 8'b00000000;
      ProductSum_for_asn_55_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_80_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_83_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_82_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_85_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_84_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_87_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_86_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_89_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_88_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_91_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_90_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_93_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_92_itm_1 <= 8'b00000000;
      ProductSum_for_asn_69_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_79_itm_1 <= 8'b00000000;
      ProductSum_for_asn_81_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_48_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_51_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_50_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_53_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_52_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_55_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_54_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_57_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_56_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_59_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_58_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_61_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_60_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_62_itm_1 <= 8'b00000000;
      ProductSum_for_asn_95_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_47_itm_1 <= 8'b00000000;
      ProductSum_for_asn_107_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_16_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_19_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_18_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_21_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_20_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_23_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_22_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_25_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_24_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_27_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_26_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_29_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_28_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_30_itm_1 <= 8'b00000000;
      ProductSum_for_asn_126_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_6_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_9_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_8_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_13_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_13_itm_1_6_0 <= 7'b0000000;
      weight_mem_run_3_for_5_mux_15_itm_1_7_6 <= 2'b00;
      weight_mem_run_3_for_5_mux_15_itm_1_5_0 <= 6'b000000;
      weight_mem_run_3_for_5_mux_14_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_14_itm_1_6_0 <= 7'b0000000;
    end
    else if ( ProductSum_for_and_cse ) begin
      ProductSum_for_asn_26_itm_6 <= ProductSum_for_asn_28_itm_5;
      ProductSum_for_asn_40_itm_6 <= ProductSum_for_asn_41_itm_5;
      weight_mem_run_3_for_5_mux_96_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_6_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_99_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_6_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_98_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_6_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      ProductSum_for_asn_55_itm_6 <= ProductSum_for_asn_56_itm_5;
      weight_mem_run_3_for_5_mux_80_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_83_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_82_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_85_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_84_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_87_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_86_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_89_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_9_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_88_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_8_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_91_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_11_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_90_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_10_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_93_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_13_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_92_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_5_12_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      ProductSum_for_asn_69_itm_6 <= ProductSum_for_asn_69_itm_5;
      weight_mem_run_3_for_5_mux_79_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_4_15_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      ProductSum_for_asn_81_itm_6 <= ProductSum_for_asn_82_itm_5;
      weight_mem_run_3_for_5_mux_48_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_51_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_50_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_53_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_52_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_55_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_54_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_57_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_9_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_56_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_8_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_59_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_11_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_58_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_10_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_61_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_13_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_60_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_12_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_62_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_14_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      ProductSum_for_asn_95_itm_6 <= ProductSum_for_asn_95_itm_5;
      weight_mem_run_3_for_5_mux_47_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_2_15_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000,
          weight_mem_run_3_for_land_3_lpi_1_dfm_2);
      ProductSum_for_asn_107_itm_6 <= ProductSum_for_asn_108_itm_5;
      weight_mem_run_3_for_5_mux_16_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_19_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_18_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_21_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_20_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_23_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_22_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_25_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_9_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_24_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_8_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_27_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_11_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_26_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_10_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_29_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_13_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_28_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_12_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_30_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_14_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      ProductSum_for_asn_126_itm_6 <= ProductSum_for_asn_128_itm_5;
      weight_mem_run_3_for_5_mux_6_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_0_6_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_9_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_0_9_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_8_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_0_8_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_13_itm_1_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_13_sva_dfm_2_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006[7]),
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_13_itm_1_6_0 <= MUX_v_7_2_2(weight_port_read_out_data_0_13_sva_dfm_2_6_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006[6:0]),
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_15_itm_1_7_6 <= MUX_v_2_2_2(weight_port_read_out_data_0_15_sva_dfm_2_7_6,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008[7:6]),
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_15_itm_1_5_0 <= MUX_v_6_2_2(weight_port_read_out_data_0_15_sva_dfm_2_5_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008[5:0]),
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_14_itm_1_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_14_sva_dfm_2_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009[7]),
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_14_itm_1_6_0 <= MUX_v_7_2_2(weight_port_read_out_data_0_14_sva_dfm_2_6_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009[6:0]),
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_214_enex5 ) begin
      weight_port_read_out_data_4_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_5_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_3 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
          <= 1'b0;
      rva_in_reg_rw_sva_6 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_cse ) begin
      weight_mem_run_3_for_land_5_lpi_1_dfm_3 <= weight_mem_run_3_for_land_5_lpi_1_dfm_2;
      weight_mem_run_3_for_land_4_lpi_1_dfm_3 <= weight_mem_run_3_for_land_4_lpi_1_dfm_2;
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= weight_mem_run_3_for_land_3_lpi_1_dfm_2;
      weight_mem_run_3_for_land_2_lpi_1_dfm_3 <= weight_mem_run_3_for_land_2_lpi_1_dfm_2;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
      rva_in_reg_rw_sva_6 <= rva_in_reg_rw_sva_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_215_enex5 ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_3_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_216_enex5 ) begin
      weight_port_read_out_data_4_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_2_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_217_enex5 ) begin
      weight_port_read_out_data_4_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_5_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_218_enex5 ) begin
      weight_port_read_out_data_4_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_4_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_219_enex5 ) begin
      weight_port_read_out_data_4_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_7_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_220_enex5 ) begin
      weight_port_read_out_data_4_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_221_enex5 ) begin
      weight_port_read_out_data_4_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_9_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_222_enex5 ) begin
      weight_port_read_out_data_4_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_8_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_223_enex5 ) begin
      weight_port_read_out_data_4_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_11_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_224_enex5 ) begin
      weight_port_read_out_data_4_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_10_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_225_enex5 ) begin
      weight_port_read_out_data_4_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_13_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_226_enex5 ) begin
      weight_port_read_out_data_4_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_12_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_227_enex5 ) begin
      weight_port_read_out_data_4_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_228_enex5 ) begin
      weight_port_read_out_data_4_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_15_enex5 ) begin
      weight_port_read_out_data_3_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_15_tmp ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
          <= MUX_v_8_2_2(8'b00000000, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_1_nl,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_229_enex5 ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_230_enex5 ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_3_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_231_enex5 ) begin
      weight_port_read_out_data_2_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_232_enex5 ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_5_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_233_enex5 ) begin
      weight_port_read_out_data_2_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_4_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_234_enex5 ) begin
      weight_port_read_out_data_2_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_7_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_235_enex5 ) begin
      weight_port_read_out_data_2_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_236_enex5 ) begin
      weight_port_read_out_data_2_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_9_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_237_enex5 ) begin
      weight_port_read_out_data_2_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_8_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_238_enex5 ) begin
      weight_port_read_out_data_2_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_11_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_239_enex5 ) begin
      weight_port_read_out_data_2_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_10_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_240_enex5 ) begin
      weight_port_read_out_data_2_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_13_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_241_enex5 ) begin
      weight_port_read_out_data_2_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_12_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_242_enex5 ) begin
      weight_port_read_out_data_2_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_243_enex5 ) begin
      weight_port_read_out_data_2_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_31_enex5 ) begin
      weight_port_read_out_data_1_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_31_tmp ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
          <= MUX_v_8_2_2(8'b00000000, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_5_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( mux_460_nl & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_0_5_sva_dfm_1_1 <= MUX1HOT_v_8_9_2(weight_port_read_out_data_0_5_sva_mx0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_cse
          , weight_mem_run_3_for_5_and_173_cse , weight_mem_run_3_for_5_and_174_cse
          , weight_mem_run_3_for_5_and_159_cse , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_177_nl , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_179_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_7_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( mux_462_nl & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_0_7_sva_dfm_1_1 <= MUX1HOT_v_8_9_2(weight_port_read_out_data_0_7_sva_mx0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_188_nl
          , weight_mem_run_3_for_5_and_173_cse , weight_mem_run_3_for_5_and_174_cse
          , weight_mem_run_3_for_5_and_191_nl , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_161_cse , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_179_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= 1'b0;
      accum_vector_operator_1_for_asn_118_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_103_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_88_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_73_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_58_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_43_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_28_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_13_itm_5 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_3_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
      accum_vector_operator_1_for_asn_118_itm_5 <= accum_vector_operator_1_for_asn_118_itm_4;
      accum_vector_operator_1_for_asn_103_itm_5 <= accum_vector_operator_1_for_asn_103_itm_4;
      accum_vector_operator_1_for_asn_88_itm_5 <= accum_vector_operator_1_for_asn_88_itm_4;
      accum_vector_operator_1_for_asn_73_itm_5 <= accum_vector_operator_1_for_asn_73_itm_4;
      accum_vector_operator_1_for_asn_58_itm_5 <= accum_vector_operator_1_for_asn_58_itm_4;
      accum_vector_operator_1_for_asn_43_itm_5 <= accum_vector_operator_1_for_asn_43_itm_4;
      accum_vector_operator_1_for_asn_28_itm_5 <= accum_vector_operator_1_for_asn_28_itm_4;
      accum_vector_operator_1_for_asn_13_itm_5 <= accum_vector_operator_1_for_asn_13_itm_4;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        & while_stage_0_6 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        & while_stage_0_6 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_5 <= 1'b0;
      rva_in_reg_rw_sva_st_5 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_3_cse ) begin
      rva_in_reg_rw_sva_st_1_5 <= rva_in_reg_rw_sva_st_1_4;
      rva_in_reg_rw_sva_st_5 <= rva_in_reg_rw_sva_st_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_2 <= 1'b0;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_28_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_30_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_31_itm_2 <= 1'b0;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= 3'b000;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2 <=
          1'b0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2 <=
          1'b0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2 <=
          1'b0;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= 3'b000;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2_cse
          <= 1'b0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse <= 1'b0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse <= 1'b0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse <= 1'b0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse <= 1'b0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_142_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_135_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_136_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_100_itm_1 <= 1'b0;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_12_itm_1 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_14_itm_1_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_16_itm_1_cse <= 1'b0;
      weight_mem_run_3_for_5_and_7_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_148_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_2 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      accum_vector_operator_1_for_asn_118_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_103_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_88_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_73_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_58_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_43_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_28_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_13_itm_4 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= 1'b0;
    end
    else if ( weight_mem_banks_read_1_read_data_and_8_cse ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_28_itm_2 <= weight_mem_run_3_for_5_and_28_itm_1;
      weight_mem_run_3_for_5_and_30_itm_2 <= weight_mem_run_3_for_5_and_30_itm_1;
      weight_mem_run_3_for_5_and_31_itm_2 <= weight_mem_run_3_for_5_and_31_itm_1;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= weight_read_addrs_7_lpi_1_dfm_2_2_0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2 <=
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_1;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2 <=
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_1;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2 <=
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_1;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= weight_read_addrs_5_lpi_1_dfm_2_2_0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2_cse
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_1;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_2_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_1;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_2_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_1;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_2_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_1;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_1;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_1;
      weight_mem_run_3_for_5_and_142_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_135_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_136_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b111)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_2_2_0!=3'b000));
      weight_mem_run_3_for_5_and_100_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b011)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
      weight_mem_run_3_for_5_and_12_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1;
      reg_weight_mem_run_3_for_5_and_14_itm_1_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1;
      reg_weight_mem_run_3_for_5_and_16_itm_1_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1;
      weight_mem_run_3_for_5_and_7_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1;
      weight_mem_run_3_for_5_and_148_itm_2 <= weight_mem_run_3_for_5_and_148_itm_1;
      weight_mem_run_3_for_5_and_150_itm_2 <= weight_mem_run_3_for_5_and_150_itm_1;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      accum_vector_operator_1_for_asn_118_itm_4 <= accum_vector_operator_1_for_asn_118_itm_3;
      accum_vector_operator_1_for_asn_103_itm_4 <= accum_vector_operator_1_for_asn_103_itm_3;
      accum_vector_operator_1_for_asn_88_itm_4 <= accum_vector_operator_1_for_asn_88_itm_3;
      accum_vector_operator_1_for_asn_73_itm_4 <= accum_vector_operator_1_for_asn_73_itm_3;
      accum_vector_operator_1_for_asn_58_itm_4 <= accum_vector_operator_1_for_asn_58_itm_3;
      accum_vector_operator_1_for_asn_43_itm_4 <= accum_vector_operator_1_for_asn_43_itm_3;
      accum_vector_operator_1_for_asn_28_itm_4 <= accum_vector_operator_1_for_asn_28_itm_3;
      accum_vector_operator_1_for_asn_13_itm_4 <= accum_vector_operator_1_for_asn_13_itm_3;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & and_dcpl_55 & weight_mem_run_3_for_land_7_lpi_1_dfm_1
        ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_18_nl) & while_stage_0_6 ) begin
      reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_28_itm_5 <= 1'b0;
      ProductSum_for_asn_41_itm_5 <= 1'b0;
      ProductSum_for_asn_56_itm_5 <= 1'b0;
      ProductSum_for_asn_82_itm_5 <= 1'b0;
      ProductSum_for_asn_108_itm_5 <= 1'b0;
      ProductSum_for_asn_128_itm_5 <= 1'b0;
      ProductSum_for_asn_69_itm_5 <= 1'b0;
      ProductSum_for_asn_95_itm_5 <= 1'b0;
    end
    else if ( ProductSum_for_and_8_cse ) begin
      ProductSum_for_asn_28_itm_5 <= ProductSum_for_asn_28_itm_4;
      ProductSum_for_asn_41_itm_5 <= ProductSum_for_asn_41_itm_4;
      ProductSum_for_asn_56_itm_5 <= ProductSum_for_asn_56_itm_4;
      ProductSum_for_asn_82_itm_5 <= ProductSum_for_asn_82_itm_4;
      ProductSum_for_asn_108_itm_5 <= ProductSum_for_asn_108_itm_4;
      ProductSum_for_asn_128_itm_5 <= ProductSum_for_asn_128_itm_4;
      ProductSum_for_asn_69_itm_5 <= ProductSum_for_asn_69_itm_4;
      ProductSum_for_asn_95_itm_5 <= ProductSum_for_asn_95_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_6_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_251) ) begin
      weight_port_read_out_data_6_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= 1'b0;
      rva_in_reg_rw_sva_5 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_4_cse ) begin
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= weight_mem_run_3_for_land_7_lpi_1_dfm_1;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1;
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= weight_mem_run_3_for_land_1_lpi_1_dfm_2;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= weight_mem_run_3_for_land_5_lpi_1_dfm_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= weight_mem_run_3_for_land_3_lpi_1_dfm_1;
      rva_in_reg_rw_sva_5 <= rva_in_reg_rw_sva_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_253) ) begin
      weight_port_read_out_data_5_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_9_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_11_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_10_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_13_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_12_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_137_cse ) begin
      weight_port_read_out_data_3_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
      weight_port_read_out_data_3_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
      weight_port_read_out_data_3_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
      weight_port_read_out_data_3_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
      weight_port_read_out_data_3_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
      weight_port_read_out_data_3_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
      weight_port_read_out_data_3_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
      weight_port_read_out_data_3_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
      weight_port_read_out_data_3_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
      weight_port_read_out_data_3_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
      weight_port_read_out_data_3_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
      weight_port_read_out_data_3_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
      weight_port_read_out_data_3_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
      weight_port_read_out_data_3_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
      weight_port_read_out_data_3_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_255) ) begin
      weight_port_read_out_data_1_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( or_939_cse & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_1_sva_dfm_1 <= weight_port_read_out_data_7_1_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_44_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_44_itm_1
          <= ~((weight_read_addrs_5_lpi_1_dfm_2_2_0!=3'b000));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_30_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2 <= 1'b0;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
          <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_375_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_30_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_30_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_1;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= weight_read_addrs_3_lpi_1_dfm_2_2_0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
          <= ~((weight_read_addrs_3_lpi_1_dfm_2_2_0!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_379_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_136_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_134_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_151_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_14_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_2
          <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_380_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_14_itm_1
          <= crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1 <= 1'b0;
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_382_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_28_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_8 <= 120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_252 | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & mux_21_nl ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_8 <= weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:8];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_252 | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)))
        ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_RunFSM_switch_lp_equal_tmp_1_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)))
        & PECore_UpdateFSM_switch_lp_equal_tmp_2_3)) & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2
          <= PECore_RunMac_PECore_RunMac_if_and_svs_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(ProductSum_for_asn_108_itm_3 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2
          <= PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_22_nl) & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_23_nl) & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ ProductSum_for_asn_41_itm_3) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_28_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1 <= 1'b0;
    end
    else if ( weight_read_addrs_and_5_cse ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_76 & (~ ProductSum_for_asn_56_itm_3) ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_76 & (~ ProductSum_for_asn_69_itm_3) ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_2_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_4_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_6_lpi_1_dfm_1_1 <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= 1'b0;
      rva_in_reg_rw_sva_4 <= 1'b0;
    end
    else if ( while_if_and_10_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_99_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_91_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_75_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp |
          Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp |
          Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 | and_749_cse
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_123_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_6_lpi_1_dfm_1_1 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & or_260_cse;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | and_747_cse
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_111_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & weight_mem_read_arbxbar_xbar_1_for_3_8_for_3_or_cse;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse;
      rva_in_reg_rw_sva_4 <= rva_in_reg_rw_sva_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_48_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_54_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_60_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_66_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_72_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_78_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_84_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_90_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva <= 15'b000000000000000;
    end
    else if ( (~ mux_464_nl) & fsm_output & while_stage_0_5 & PECoreRun_wen ) begin
      pe_manager_base_weight_sva <= pe_manager_base_weight_sva_mx2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= 11'b00000000000;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= 1'b0;
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_371_itm_1 <= 1'b0;
      rva_in_reg_rw_sva_3 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= 1'b0;
    end
    else if ( weight_read_addrs_and_7_cse ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= MUX_v_11_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl,
          weight_read_addrs_0_14_4_lpi_1_dfm_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= MUX_s_1_2_2((weight_read_addrs_0_3_0_lpi_1_dfm_4[3]),
          (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= nor_375_cse;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1 <= MUX_s_1_2_2((pe_manager_base_weight_sva_mx1_3_0[2]),
          reg_rva_in_reg_rw_sva_2_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_371_itm_1 <= MUX_s_1_2_2(pe_manager_base_weight_sva_mx3_0,
          reg_rva_in_reg_rw_sva_2_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      rva_in_reg_rw_sva_3 <= reg_rva_in_reg_rw_sva_2_cse;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_155 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_48_enex5 ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_15_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_49_enex5 ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_14_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_50_enex5 ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_13_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_51_enex5 ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_12_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_52_enex5 ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_11_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_53_enex5 ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_10_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_54_enex5 ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_9_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_55_enex5 ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_8_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_56_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_57_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_58_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_59_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_60_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_61_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_62_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_63_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= 12'b000000000000;
    end
    else if ( weight_write_addrs_and_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= weight_write_addrs_lpi_1_dfm_1_2[14:3];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= 1'b0;
      weight_read_addrs_1_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_3_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= 13'b0000000000000;
      weight_read_addrs_5_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_7_lpi_1_dfm_1 <= 15'b000000000000000;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= 1'b0;
      accum_vector_operator_1_for_asn_118_itm_2 <= 1'b0;
      accum_vector_operator_1_for_asn_103_itm_2 <= 1'b0;
      accum_vector_operator_1_for_asn_88_itm_2 <= 1'b0;
      accum_vector_operator_1_for_asn_58_itm_2 <= 1'b0;
      accum_vector_operator_1_for_asn_13_itm_2 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1,
          and_156_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1,
          and_156_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1,
          and_156_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1,
          and_156_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1,
          and_156_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1,
          and_156_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1,
          and_156_cse);
      weight_read_addrs_1_lpi_1_dfm_1 <= weight_read_addrs_1_lpi_1_dfm_1_1;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_3_lpi_1_dfm_1 <= weight_read_addrs_3_lpi_1_dfm_1_1;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_1 <= weight_read_addrs_5_lpi_1_dfm_1_1;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_7_lpi_1_dfm_1 <= weight_read_addrs_7_lpi_1_dfm_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_34_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_tmp;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_not_185,
          weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0, and_107_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0, and_114_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0, and_121_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0, and_dcpl_598);
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0, and_135_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0, and_142_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0, and_dcpl_619);
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0, and_156_cse);
      accum_vector_operator_1_for_asn_118_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2;
      accum_vector_operator_1_for_asn_103_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2;
      accum_vector_operator_1_for_asn_88_itm_2 <= accum_vector_operator_1_for_asn_88_itm_1;
      accum_vector_operator_1_for_asn_58_itm_2 <= PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2;
      accum_vector_operator_1_for_asn_13_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_25_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= 8'b00000000;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_15_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_requests_transpose_and_13_cse ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= weight_mem_write_arbxbar_xbar_for_lshift_tmp;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_15_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b101)
          & nor_375_cse;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b011)
          & nor_375_cse;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b110)
          & nor_375_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_and_cse ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_576);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_576);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_576);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_576);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_576);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_576);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_576);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_576);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_64_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( weight_read_addrs_and_7_cse & ((~ while_stage_0_5) | while_and_1263_itm_1)
        ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= MUX_v_15_2_2(pe_manager_base_weight_sva_mx2,
          PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1, while_and_1263_itm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_64_enex5 ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_15_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_65_enex5 ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_14_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_66_enex5 ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_13_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_67_enex5 ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_12_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_68_enex5 ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_11_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_69_enex5 ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_10_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_70_enex5 ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_9_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_71_enex5 ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_8_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_72_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_7_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_73_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_6_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_74_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_5_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_75_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_76_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_3_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_77_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_2_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_78_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_1_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_79_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= 15'b000000000000000;
    end
    else if ( weight_write_addrs_and_2_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= pe_manager_base_input_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= 1'b0;
      reg_rva_in_reg_rw_sva_2_cse <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= 1'b0;
      while_and_1263_itm_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiWrite_switch_lp_and_2_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(accum_vector_data_3_sva_1_load_mx0w1,
          PECore_DecodeAxiWrite_switch_lp_equal_tmp_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      reg_rva_in_reg_rw_sva_2_cse <= reg_rva_in_reg_rw_sva_st_1_1_cse;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= MUX_s_1_2_2(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
      while_and_1263_itm_1 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1
          & PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
          & reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= 4'b0000;
    end
    else if ( weight_read_addrs_and_29_enex5 ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= 11'b00000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_209 ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_2_1_sva <= 2'b00;
      pe_config_is_zero_first_sva <= 1'b0;
    end
    else if ( state_and_cse ) begin
      state_2_1_sva <= state_mux_1_cse;
      pe_config_is_zero_first_sva <= pe_config_is_zero_first_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_0_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_259) ) begin
      state_0_sva <= PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_manager_counter_sva <= 4'b0000;
    end
    else if ( (((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4:2]!=3'b000))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:5]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10:8]!=3'b000))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:11]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
        & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])
        & rva_in_PopNB_mioi_return_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]==2'b00)
        & and_dcpl_214) | and_1287_cse) & PECoreRun_wen ) begin
      pe_config_manager_counter_sva <= MUX_v_4_2_2(pe_config_manager_counter_sva_dfm_3_1,
          PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl,
          and_638_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_num_manager_sva <= 4'b0001;
      pe_config_num_output_sva <= 8'b00000001;
    end
    else if ( pe_config_num_manager_and_cse ) begin
      pe_config_num_manager_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[35:32];
      pe_config_num_output_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= 1'b0;
      state_2_1_sva_dfm_1 <= 2'b00;
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= 8'b00000000;
      input_write_req_valid_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_5_cse ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= rva_in_PopNB_mioi_return_rsc_z_mxwt;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
      state_2_1_sva_dfm_1 <= MUX_v_2_2_2(PECore_UpdateFSM_switch_lp_and_1_nl, state_mux_1_cse,
          rva_in_PopNB_mioi_return_rsc_z_mxwt);
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= and_315_cse;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0];
      input_write_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= 1'b0;
      PECore_RunFSM_switch_lp_nor_tmp_1 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_9_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= PECore_UpdateFSM_switch_lp_equal_tmp_6;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= ~(PECore_RunScale_PECore_RunScale_if_and_1_svs_1
          | PECore_UpdateFSM_switch_lp_nor_tmp_1);
      PECore_RunFSM_switch_lp_nor_tmp_1 <= ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
          | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(or_407_cse | or_dcpl_259)) ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= input_port_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva <= 8'b00000000;
    end
    else if ( or_945_cse & mux_465_nl & and_dcpl_949 & PECoreRun_wen ) begin
      pe_config_input_counter_sva <= pe_config_input_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva <= 8'b00000000;
    end
    else if ( or_945_cse & mux_466_nl & and_dcpl_949 & PECoreRun_wen ) begin
      pe_config_output_counter_sva <= pe_config_output_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      operator_8_false_acc_sdt_sva_1 <= 9'b000000000;
    end
    else if ( pe_config_UpdateManagerCounter_if_if_and_enex5 ) begin
      operator_8_false_acc_sdt_sva_1 <= nl_operator_8_false_acc_sdt_sva_1[8:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiWrite_switch_lp_and_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_244_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd <= weight_port_read_out_data_0_1_sva_dfm_2_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_245_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1 <= weight_port_read_out_data_0_1_sva_dfm_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd <= 1'b0;
      reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_138_cse ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd <= weight_port_read_out_data_0_2_sva_dfm_2_rsp_0;
      reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd <= weight_port_read_out_data_0_3_sva_dfm_2_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_246_enex5 ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_1 <= weight_port_read_out_data_0_2_sva_dfm_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_1_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[15:8]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_189_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_199_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_202_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[23:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_203_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_2_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[15:8]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_219_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_229_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_230_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_232_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= 1'b0;
    end
    else if ( weight_read_addrs_and_17_cse ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= 1'b0;
    end
    else if ( PECoreRun_wen & weight_mem_run_3_for_land_5_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2 <= 2'b00;
    end
    else if ( PECoreRun_wen & mux_35_nl & while_stage_0_6 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2 <= MUX_v_2_2_2(pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_2[7:6]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_9_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_11_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_10_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_13_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_12_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_15_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_143_cse ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_9_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_11_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_10_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_13_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_12_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_158_cse ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
      weight_port_read_out_data_5_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
      weight_port_read_out_data_5_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
      weight_port_read_out_data_5_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
      weight_port_read_out_data_5_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
      weight_port_read_out_data_5_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
      weight_port_read_out_data_5_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
      weight_port_read_out_data_5_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
      weight_port_read_out_data_5_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
      weight_port_read_out_data_5_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
      weight_port_read_out_data_5_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
      weight_port_read_out_data_5_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
      weight_port_read_out_data_5_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_run_3_for_land_5_lpi_1_dfm_2) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
        | (~ while_stage_0_7))) ) begin
      weight_port_read_out_data_4_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_run_3_for_land_3_lpi_1_dfm_2) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
        | (~ while_stage_0_7))) ) begin
      weight_port_read_out_data_2_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_9_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_11_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_10_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_13_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_12_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_185_cse ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
      weight_port_read_out_data_1_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
      weight_port_read_out_data_1_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
      weight_port_read_out_data_1_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
      weight_port_read_out_data_1_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
      weight_port_read_out_data_1_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
      weight_port_read_out_data_1_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
      weight_port_read_out_data_1_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
      weight_port_read_out_data_1_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
      weight_port_read_out_data_1_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
      weight_port_read_out_data_1_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
      weight_port_read_out_data_1_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
      weight_port_read_out_data_1_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
      weight_port_read_out_data_1_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_6_sva_dfm_2 <= 8'b00000000;
      weight_port_read_out_data_0_9_sva_dfm_2 <= 8'b00000000;
      weight_port_read_out_data_0_8_sva_dfm_2 <= 8'b00000000;
      weight_port_read_out_data_0_11_sva_dfm_2 <= 8'b00000000;
      weight_port_read_out_data_0_12_sva_dfm_2 <= 8'b00000000;
      weight_port_read_out_data_0_13_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_13_sva_dfm_2_6_0 <= 7'b0000000;
      weight_port_read_out_data_0_15_sva_dfm_2_7_6 <= 2'b00;
      weight_port_read_out_data_0_15_sva_dfm_2_5_0 <= 6'b000000;
      weight_port_read_out_data_0_14_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_14_sva_dfm_2_6_0 <= 7'b0000000;
      weight_port_read_out_data_0_10_sva_dfm_2_7_4 <= 4'b0000;
      weight_port_read_out_data_0_10_sva_dfm_2_3_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_199_cse ) begin
      weight_port_read_out_data_0_6_sva_dfm_2 <= MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_sva_1,
          while_and_40_tmp);
      weight_port_read_out_data_0_9_sva_dfm_2 <= MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_sva_1,
          while_and_40_tmp);
      weight_port_read_out_data_0_8_sva_dfm_2 <= MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_sva_1,
          while_and_40_tmp);
      weight_port_read_out_data_0_11_sva_dfm_2 <= MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1,
          while_and_40_tmp);
      weight_port_read_out_data_0_12_sva_dfm_2 <= MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_sva_1,
          while_and_40_tmp);
      weight_port_read_out_data_0_13_sva_dfm_2_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006[7]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000,
          while_and_40_tmp);
      weight_port_read_out_data_0_13_sva_dfm_2_6_0 <= MUX_v_7_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006[6:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001,
          while_and_40_tmp);
      weight_port_read_out_data_0_15_sva_dfm_2_7_6 <= MUX_v_2_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008[7:6]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000,
          while_and_40_tmp);
      weight_port_read_out_data_0_15_sva_dfm_2_5_0 <= MUX_v_6_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008[5:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000001,
          while_and_40_tmp);
      weight_port_read_out_data_0_14_sva_dfm_2_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009[7]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000,
          while_and_40_tmp);
      weight_port_read_out_data_0_14_sva_dfm_2_6_0 <= MUX_v_7_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009[6:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001,
          while_and_40_tmp);
      weight_port_read_out_data_0_10_sva_dfm_2_7_4 <= MUX_v_4_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005[7:4]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000000,
          while_and_40_tmp);
      weight_port_read_out_data_0_10_sva_dfm_2_3_0 <= MUX_v_4_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005[3:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000001,
          while_and_40_tmp);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_15_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1279_cse | or_dcpl_390 | weight_mem_run_3_for_5_and_28_itm_2)
        & and_dcpl_958 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_15_sva_dfm_1_1 <= weight_port_read_out_data_7_15_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_14_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1327_cse | or_dcpl_395 | or_dcpl_394) & and_dcpl_958 & PECoreRun_wen
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_14_sva_dfm_1_1 <= weight_port_read_out_data_7_14_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_13_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1332_cse | weight_mem_run_3_for_5_and_135_itm_1 | weight_mem_run_3_for_5_and_142_itm_1
        | weight_mem_run_3_for_5_and_28_itm_2) & and_dcpl_958 & PECoreRun_wen & (~
        while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_13_sva_dfm_1_1 <= weight_port_read_out_data_7_13_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_12_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1332_cse | or_dcpl_403 | weight_mem_run_3_for_5_and_28_itm_2)
        & and_dcpl_958 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_12_sva_dfm_1_1 <= weight_port_read_out_data_7_12_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_11_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1327_cse | or_dcpl_408 | or_dcpl_407) & and_dcpl_958 & PECoreRun_wen
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_11_sva_dfm_1_1 <= weight_port_read_out_data_7_11_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_10_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1327_cse | or_dcpl_395 | weight_mem_run_3_for_5_and_30_itm_2 |
        weight_mem_run_3_for_5_and_100_itm_1) & and_dcpl_958 & PECoreRun_wen & (~
        while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_10_sva_dfm_1_1 <= weight_port_read_out_data_7_10_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_9_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1352_cse | or_dcpl_395 | or_dcpl_407) & and_dcpl_958 & PECoreRun_wen
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_9_sva_dfm_1_1 <= weight_port_read_out_data_7_9_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_8_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( or_939_cse & and_dcpl_958 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_8_sva_dfm_1_1 <= weight_port_read_out_data_7_8_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_7_sva_dfm_1_1 <= 8'b00000000;
      weight_port_read_out_data_7_6_sva_dfm_1_1 <= 8'b00000000;
      weight_port_read_out_data_7_5_sva_dfm_1_1 <= 8'b00000000;
      weight_port_read_out_data_7_4_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( and_1363_cse ) begin
      weight_port_read_out_data_7_7_sva_dfm_1_1 <= weight_port_read_out_data_7_7_sva_dfm_1_2;
      weight_port_read_out_data_7_6_sva_dfm_1_1 <= weight_port_read_out_data_7_6_sva_dfm_1_2;
      weight_port_read_out_data_7_5_sva_dfm_1_1 <= weight_port_read_out_data_7_5_sva_dfm_1_2;
      weight_port_read_out_data_7_4_sva_dfm_1_1 <= weight_port_read_out_data_7_4_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_3_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1332_cse | or_dcpl_403 | weight_mem_run_3_for_5_and_100_itm_1)
        & and_dcpl_958 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_3_sva_dfm_1_1 <= weight_port_read_out_data_7_3_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_2_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1332_cse | or_dcpl_390 | weight_mem_run_3_for_5_and_100_itm_1)
        & and_dcpl_958 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_2_sva_dfm_1_1 <= weight_port_read_out_data_7_2_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_0_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1352_cse | or_dcpl_395 | weight_mem_run_3_for_5_and_142_itm_1
        | weight_mem_run_3_for_5_and_100_itm_1) & and_dcpl_958 & PECoreRun_wen &
        (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_0_sva_dfm_1_1 <= weight_port_read_out_data_7_0_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_15_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1397_cse | reg_weight_mem_run_3_for_5_and_16_itm_1_cse | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_2_cse_2
        | reg_weight_mem_run_3_for_5_and_14_itm_1_cse | weight_mem_run_3_for_5_and_12_itm_1)
        & and_dcpl_958 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_5_15_sva_dfm_1_1 <= weight_port_read_out_data_5_15_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_14_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1397_cse | reg_weight_mem_run_3_for_5_and_16_itm_1_cse | weight_mem_run_3_for_5_and_7_itm_1
        | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_2_cse_2
        | reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_2_cse_2)
        & and_dcpl_958 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_5_14_sva_dfm_1_1 <= weight_port_read_out_data_5_14_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_384_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
          <= MUX_s_1_2_2(weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_1,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_36_nl & while_stage_0_6 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= 8'b00000000;
    end
    else if ( mux_490_nl & and_dcpl_958 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_37_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= MUX_v_8_2_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[7:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_48_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_38_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= MUX_v_8_2_2((weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[7:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_80_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_5_and_31_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_30_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_28_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_1
          <= 1'b0;
      weight_mem_run_3_for_land_lpi_1_dfm_1_1 <= 1'b0;
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_148_itm_1 <= 1'b0;
      accum_vector_operator_1_for_asn_118_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_103_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_88_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_73_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_58_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_43_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_28_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_13_itm_3 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= 1'b0;
    end
    else if ( weight_read_addrs_and_19_cse ) begin
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= weight_read_addrs_5_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_5_and_31_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_30_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_28_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_1[2:0]!=3'b000));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_359_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_358_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_356_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_121_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_119_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_1
          <= ~((pe_manager_base_weight_sva[2:0]!=3'b000));
      weight_mem_run_3_for_land_lpi_1_dfm_1_1 <= weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= weight_read_addrs_7_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= ~((weight_read_addrs_5_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_150_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1
          & (pe_manager_base_weight_sva[1:0]==2'b01) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_148_itm_1 <= (pe_manager_base_weight_sva[1]) & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_371_itm_1
          & (~ (pe_manager_base_weight_sva[2])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      accum_vector_operator_1_for_asn_118_itm_3 <= accum_vector_operator_1_for_asn_118_itm_2;
      accum_vector_operator_1_for_asn_103_itm_3 <= accum_vector_operator_1_for_asn_103_itm_2;
      accum_vector_operator_1_for_asn_88_itm_3 <= accum_vector_operator_1_for_asn_88_itm_2;
      accum_vector_operator_1_for_asn_73_itm_3 <= accum_vector_operator_1_for_asn_73_itm_2;
      accum_vector_operator_1_for_asn_58_itm_3 <= accum_vector_operator_1_for_asn_58_itm_2;
      accum_vector_operator_1_for_asn_43_itm_3 <= accum_vector_operator_1_for_asn_43_itm_2;
      accum_vector_operator_1_for_asn_28_itm_3 <= accum_vector_operator_1_for_asn_28_itm_2;
      accum_vector_operator_1_for_asn_13_itm_3 <= accum_vector_operator_1_for_asn_13_itm_2;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_30_itm_1
          <= 1'b0;
    end
    else if ( weight_read_addrs_and_20_cse ) begin
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= weight_read_addrs_3_lpi_1_dfm_1[2:0];
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_30_itm_1
          <= ~((weight_read_addrs_3_lpi_1_dfm_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        | (~ while_stage_0_6))) ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        | (~ while_stage_0_6))) ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        | (~ while_stage_0_6))) ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_43_nl ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_60_nl ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_62_nl ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_30_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= 1'b0;
    end
    else if ( operator_15_false_1_and_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_156_cse | or_237_cse)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_dcpl_619 | or_237_cse)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_142_cse | or_237_cse)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_135_cse | or_237_cse)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_dcpl_598 | or_237_cse)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_121_cse | or_237_cse)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_114_cse | or_237_cse)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= 15'b000000000000000;
    end
    else if ( PEManager_15U_PEManagerWrite_and_enex5 ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= rva_in_reg_data_sva_1[30:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_num_input_sva <= 8'b00000001;
      pe_manager_base_bias_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_num_input_and_cse ) begin
      pe_manager_num_input_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      pe_manager_base_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[46:32];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_is_valid_sva <= 1'b0;
      pe_config_is_cluster_sva <= 1'b0;
      pe_config_is_bias_sva <= 1'b0;
    end
    else if ( pe_config_is_valid_and_cse ) begin
      pe_config_is_valid_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
      pe_config_is_cluster_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[16];
      pe_config_is_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_zero_active_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & and_315_cse & (~ PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)
        & (~ or_dcpl_270) ) begin
      pe_manager_zero_active_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:2]==8'b00000000) & nor_589_cse
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:12]!=2'b00))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:14]!=2'b00)))
        & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]))
        | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
        | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 | (~(reg_rva_in_reg_rw_sva_st_1_1_cse
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
        & while_stage_0_3))) & rva_in_PopNB_mioi_return_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100)
        & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & rva_in_reg_rw_and_5_cse ) begin
      pe_config_output_counter_sva_dfm_1 <= MUX_v_8_2_2(8'b00000000, pe_config_output_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1434_tmp ) begin
      pe_config_input_counter_sva_dfm_1 <= MUX_v_8_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl,
          PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_1_nl,
          rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_mux_27_itm_1 <= 1'b0;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= 4'b0000;
      weight_write_data_data_0_15_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_14_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_13_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_12_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_11_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_10_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_9_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_8_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= 11'b00000000000;
    end
    else if ( while_if_and_14_cse ) begin
      while_if_mux_27_itm_1 <= MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_27_nl,
          rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:0])
          & ({{3{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_4_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
      weight_write_data_data_0_15_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:120])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_14_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[119:112])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_13_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:104])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_12_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[103:96])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_11_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:88])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_10_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[87:80])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_9_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:72])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_8_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:4])
          & ({{10{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_11_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= 1'b0;
    end
    else if ( PECoreRun_wen & (and_dcpl_29 | and_dcpl_277) ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & not_tmp_33 & while_stage_0_7 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_4 <= 1'b0;
      rva_in_reg_rw_sva_st_4 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_6_cse ) begin
      rva_in_reg_rw_sva_st_1_4 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_371_itm_1;
      rva_in_reg_rw_sva_st_4 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_7 <= 1'b0;
      rva_in_reg_rw_sva_st_7 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_7_cse ) begin
      rva_in_reg_rw_sva_st_1_7 <= rva_in_reg_rw_sva_st_1_6;
      rva_in_reg_rw_sva_st_7 <= rva_in_reg_rw_sva_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= 4'b0000;
    end
    else if ( PECoreRun_wen & and_dcpl_263 ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_28_itm_4 <= 1'b0;
      ProductSum_for_asn_41_itm_4 <= 1'b0;
      ProductSum_for_asn_56_itm_4 <= 1'b0;
      ProductSum_for_asn_82_itm_4 <= 1'b0;
      ProductSum_for_asn_108_itm_4 <= 1'b0;
      ProductSum_for_asn_128_itm_4 <= 1'b0;
      ProductSum_for_asn_69_itm_4 <= 1'b0;
      ProductSum_for_asn_95_itm_4 <= 1'b0;
    end
    else if ( ProductSum_for_and_14_cse ) begin
      ProductSum_for_asn_28_itm_4 <= ProductSum_for_asn_28_itm_3;
      ProductSum_for_asn_41_itm_4 <= ProductSum_for_asn_41_itm_3;
      ProductSum_for_asn_56_itm_4 <= ProductSum_for_asn_56_itm_3;
      ProductSum_for_asn_82_itm_4 <= ProductSum_for_asn_82_itm_3;
      ProductSum_for_asn_108_itm_4 <= ProductSum_for_asn_108_itm_3;
      ProductSum_for_asn_128_itm_4 <= ProductSum_for_asn_128_itm_3;
      ProductSum_for_asn_69_itm_4 <= ProductSum_for_asn_69_itm_3;
      ProductSum_for_asn_95_itm_4 <= ProductSum_for_asn_95_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_404_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_135_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_142_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_132_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_408_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_15_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= MUX_v_3_2_2((weight_read_addrs_1_lpi_1_dfm_1[2:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2
          <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_152_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b101)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b011)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_1 <= (pe_manager_base_weight_sva[2])
          & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_1 <= (pe_manager_base_weight_sva[1])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 & (~
          (pe_manager_base_weight_sva[2])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1
          <= ~((pe_manager_base_weight_sva[2:1]!=2'b00) | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1 <= (pe_manager_base_weight_sva[2])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1 & (pe_manager_base_weight_sva[0])
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1
          & (pe_manager_base_weight_sva[1:0]==2'b10) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1 <= (pe_manager_base_weight_sva[2])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 & (~
          (pe_manager_base_weight_sva[1])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 & (~
          (pe_manager_base_weight_sva[1])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1
          <= ~(pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1 |
          (pe_manager_base_weight_sva[1:0]!=2'b00));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1
          & (pe_manager_base_weight_sva[0]) & (~ (pe_manager_base_weight_sva[2]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_9_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_39_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_40_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_41_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_42_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_6_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_8 <= 1'b0;
    end
    else if ( PECoreRun_wen & (and_dcpl_284 | and_dcpl_277) ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_8 <= PECore_RunMac_PECore_RunMac_if_and_svs_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & or_260_cse & and_dcpl_248 ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_30_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= 1'b0;
      reg_rva_out_reg_data_127_120_sva_dfm_4_3_ftd <= 2'b00;
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd <= 1'b0;
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( input_read_req_valid_and_1_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= input_read_req_valid_lpi_1_dfm_1_7;
      reg_rva_out_reg_data_127_120_sva_dfm_4_3_ftd <= rva_out_reg_data_127_120_sva_dfm_4_2_rsp_0;
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd <= rva_out_reg_data_119_112_sva_dfm_4_2_rsp_0;
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd <= rva_out_reg_data_111_104_sva_dfm_4_2_rsp_0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_7_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_6_1 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_143_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_6_1 <= rva_out_reg_data_30_25_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_6 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_144_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_6 <= rva_out_reg_data_23_17_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_145_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= rva_out_reg_data_15_9_sva_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_247_enex5 ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd_1 <= weight_port_read_out_data_0_3_sva_dfm_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_146_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= rva_out_reg_data_35_32_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_147_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_3 <= rva_out_reg_data_39_36_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_148_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3 <= rva_out_reg_data_46_40_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_149_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_3 <= rva_out_reg_data_62_56_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_150_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3 <= rva_out_reg_data_55_48_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_3_ftd_1 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_151_enex5 ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_3_ftd_1 <= rva_out_reg_data_127_120_sva_dfm_4_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_152_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd_1 <= rva_out_reg_data_119_112_sva_dfm_4_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_153_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd_1 <= rva_out_reg_data_111_104_sva_dfm_4_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_88_sva_dfm_4_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_154_enex5 ) begin
      rva_out_reg_data_95_88_sva_dfm_4_3 <= rva_out_reg_data_95_88_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_72_sva_dfm_4_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_155_enex5 ) begin
      rva_out_reg_data_79_72_sva_dfm_4_3 <= rva_out_reg_data_79_72_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_4_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_156_enex5 ) begin
      rva_out_reg_data_71_64_sva_dfm_4_3 <= rva_out_reg_data_71_64_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_284 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_4_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_250_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_175_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_190_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_205_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_220_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_251_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_176_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_191_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_206_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_221_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_252_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_177_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_192_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_207_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_222_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_253_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_178_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_193_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_208_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_223_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_254_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_179_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_194_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_209_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_224_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_255_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_180_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_195_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_210_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_225_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_241_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_181_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_196_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_211_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_226_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_242_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_257_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_182_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_197_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_212_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_227_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_243_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_183_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_198_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_213_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_228_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1
          <= 8'b00000000;
    end
    else if ( mux_497_nl & PECoreRun_wen ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1
          <= MUX_v_8_2_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_nl,
          weight_port_read_out_data_0_7_sva_dfm_mx0w1, or_dcpl_249);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1
          <= 8'b00000000;
    end
    else if ( mux_503_nl & PECoreRun_wen ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1
          <= MUX_v_8_2_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_nl,
          weight_port_read_out_data_0_5_sva_dfm_mx0w1, or_dcpl_249);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_56_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_244_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_245_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_247_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[23:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_248_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_57_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= MUX_v_8_2_2(8'b00000000, mux1h_6_nl, not_2283_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= MUX_v_8_2_2(8'b00000000, mux1h_7_nl, not_2285_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1
          <= MUX_v_8_2_2(8'b00000000, mux1h_8_nl, not_2287_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_62_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_200_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_201_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_64_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_246_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[7:0]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_140_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_67_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_231_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[23:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_233_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= 8'b00000000;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_empty_and_enex5 ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= weight_mem_write_arbxbar_xbar_for_empty_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_data_sva_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rva_in_reg_data_and_tmp ) begin
      rva_in_reg_data_sva_1 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & nand_41_cse & while_stage_0_8 ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
        & while_stage_0_6 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]))) & while_stage_0_4 )
        begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_6 <= 1'b0;
      rva_in_reg_rw_sva_st_6 <= 1'b0;
      PECore_PushAxiRsp_mux_23_itm_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_10_cse ) begin
      rva_in_reg_rw_sva_st_1_6 <= rva_in_reg_rw_sva_st_1_5;
      rva_in_reg_rw_sva_st_6 <= rva_in_reg_rw_sva_st_5;
      PECore_PushAxiRsp_mux_23_itm_1 <= MUX_s_1_2_2(weight_port_read_out_data_mux_106_nl,
          rva_out_reg_data_63_sva_dfm_7, rva_in_reg_rw_sva_5);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_28_itm_3 <= 1'b0;
      ProductSum_for_asn_41_itm_3 <= 1'b0;
      ProductSum_for_asn_56_itm_3 <= 1'b0;
      ProductSum_for_asn_108_itm_3 <= 1'b0;
      ProductSum_for_asn_128_itm_3 <= 1'b0;
      ProductSum_for_asn_69_itm_3 <= 1'b0;
    end
    else if ( ProductSum_for_and_22_cse ) begin
      ProductSum_for_asn_28_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_28_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_41_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_41_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_56_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_56_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_108_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_108_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_128_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_128_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_69_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_69_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_82_itm_3 <= 1'b0;
      ProductSum_for_asn_95_itm_3 <= 1'b0;
    end
    else if ( ProductSum_for_and_26_cse ) begin
      ProductSum_for_asn_82_itm_3 <= ProductSum_for_asn_82_itm_2;
      ProductSum_for_asn_95_itm_3 <= ProductSum_for_asn_95_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_410_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_1 <= 2'b00;
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= 1'b0;
    end
    else if ( pe_manager_base_weight_and_5_cse ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_1 <= pe_manager_base_weight_sva[1:0];
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= weight_read_addrs_4_14_2_lpi_1_dfm_1[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_1 <= 1'b0;
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( pe_manager_base_weight_and_6_cse ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_1 <= pe_manager_base_weight_sva[0];
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse
        & and_dcpl_248 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_1
          <= ~((weight_read_addrs_1_lpi_1_dfm_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_158_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1,
          ProductSum_for_asn_69_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1,
          ProductSum_for_asn_56_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          ProductSum_for_asn_41_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          ProductSum_for_asn_28_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          ProductSum_for_asn_128_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1,
          PECore_UpdateFSM_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1,
          PECore_RunFSM_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1,
          ProductSum_for_asn_108_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_73_nl & while_stage_0_5 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          accum_vector_operator_1_for_asn_73_itm_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_18_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_43_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= weight_mem_run_3_for_5_mux_11_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_44_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= weight_mem_run_3_for_5_mux_107_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_45_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= weight_mem_run_3_for_5_mux_108_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_46_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= weight_mem_run_3_for_5_mux_109_itm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_7_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_74_nl & while_stage_0_8 ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_7 <= PECore_RunMac_PECore_RunMac_if_and_svs_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= 1'b0;
      rva_out_reg_data_127_120_sva_dfm_4_2_rsp_0 <= 2'b00;
      rva_out_reg_data_119_112_sva_dfm_4_2_rsp_0 <= 1'b0;
      rva_out_reg_data_111_104_sva_dfm_4_2_rsp_0 <= 1'b0;
    end
    else if ( input_read_req_valid_and_2_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= input_read_req_valid_lpi_1_dfm_1_6;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
      rva_out_reg_data_127_120_sva_dfm_4_2_rsp_0 <= rva_out_reg_data_127_120_sva_dfm_4_1_7_6;
      rva_out_reg_data_119_112_sva_dfm_4_2_rsp_0 <= rva_out_reg_data_119_112_sva_dfm_4_1_7;
      rva_out_reg_data_111_104_sva_dfm_4_2_rsp_0 <= rva_out_reg_data_111_104_sva_dfm_4_1_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_11_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_157_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= weight_mem_run_3_for_5_mux_12_itm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_158_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= weight_mem_run_3_for_5_mux_111_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_7 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_159_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_7 <= weight_mem_run_3_for_5_mux_110_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_160_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= rva_out_reg_data_35_32_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_161_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_2 <= rva_out_reg_data_39_36_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_162_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2 <= rva_out_reg_data_46_40_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_163_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_2 <= rva_out_reg_data_62_56_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_164_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2 <= rva_out_reg_data_55_48_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_88_sva_dfm_4_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_165_enex5 ) begin
      rva_out_reg_data_95_88_sva_dfm_4_2 <= rva_out_reg_data_95_88_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_72_sva_dfm_4_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_166_enex5 ) begin
      rva_out_reg_data_79_72_sva_dfm_4_2 <= rva_out_reg_data_79_72_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_4_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_167_enex5 ) begin
      rva_out_reg_data_71_64_sva_dfm_4_2 <= rva_out_reg_data_71_64_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_33 & ((~ PECore_UpdateFSM_switch_lp_equal_tmp_2_6)
        | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6) ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
        & rva_in_reg_rw_sva_st_1_5)) & while_stage_0_7 ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5,
          (weight_port_read_out_data_0_5_sva_dfm_mx0w1[7]), PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_40_tmp , while_and_39_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= 1'b0;
      accum_vector_operator_1_for_asn_88_itm_1 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_8_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
      accum_vector_operator_1_for_asn_88_itm_1 <= accum_vector_data_5_sva_1_load_mx0w0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_28_itm_2 <= 1'b0;
      ProductSum_for_asn_41_itm_2 <= 1'b0;
      ProductSum_for_asn_56_itm_2 <= 1'b0;
      ProductSum_for_asn_82_itm_2 <= 1'b0;
      ProductSum_for_asn_108_itm_2 <= 1'b0;
      ProductSum_for_asn_128_itm_2 <= 1'b0;
      ProductSum_for_asn_69_itm_2 <= 1'b0;
      ProductSum_for_asn_95_itm_2 <= 1'b0;
    end
    else if ( ProductSum_for_and_30_cse ) begin
      ProductSum_for_asn_28_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
      ProductSum_for_asn_41_itm_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
      ProductSum_for_asn_56_itm_2 <= ProductSum_for_asn_56_itm_1;
      ProductSum_for_asn_82_itm_2 <= ProductSum_for_asn_82_itm_1;
      ProductSum_for_asn_108_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1;
      ProductSum_for_asn_128_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
      ProductSum_for_asn_69_itm_2 <= ProductSum_for_asn_69_itm_1;
      ProductSum_for_asn_95_itm_2 <= ProductSum_for_asn_95_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_27_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_4[0];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_4[8];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[16];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[31];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= MUX_v_128_256_2(input_mem_banks_bank_a_0_sva_dfm_2,
          input_mem_banks_bank_a_1_sva_dfm_2, input_mem_banks_bank_a_2_sva_dfm_2,
          input_mem_banks_bank_a_3_sva_dfm_2, input_mem_banks_bank_a_4_sva_dfm_2,
          input_mem_banks_bank_a_5_sva_dfm_2, input_mem_banks_bank_a_6_sva_dfm_2,
          input_mem_banks_bank_a_7_sva_dfm_2, input_mem_banks_bank_a_8_sva_dfm_2,
          input_mem_banks_bank_a_9_sva_dfm_2, input_mem_banks_bank_a_10_sva_dfm_2,
          input_mem_banks_bank_a_11_sva_dfm_2, input_mem_banks_bank_a_12_sva_dfm_2,
          input_mem_banks_bank_a_13_sva_dfm_2, input_mem_banks_bank_a_14_sva_dfm_2,
          input_mem_banks_bank_a_15_sva_dfm_2, input_mem_banks_bank_a_16_sva_dfm_2,
          input_mem_banks_bank_a_17_sva_dfm_2, input_mem_banks_bank_a_18_sva_dfm_2,
          input_mem_banks_bank_a_19_sva_dfm_2, input_mem_banks_bank_a_20_sva_dfm_2,
          input_mem_banks_bank_a_21_sva_dfm_2, input_mem_banks_bank_a_22_sva_dfm_2,
          input_mem_banks_bank_a_23_sva_dfm_2, input_mem_banks_bank_a_24_sva_dfm_2,
          input_mem_banks_bank_a_25_sva_dfm_2, input_mem_banks_bank_a_26_sva_dfm_2,
          input_mem_banks_bank_a_27_sva_dfm_2, input_mem_banks_bank_a_28_sva_dfm_2,
          input_mem_banks_bank_a_29_sva_dfm_2, input_mem_banks_bank_a_30_sva_dfm_2,
          input_mem_banks_bank_a_31_sva_dfm_2, input_mem_banks_bank_a_32_sva_dfm_2,
          input_mem_banks_bank_a_33_sva_dfm_2, input_mem_banks_bank_a_34_sva_dfm_2,
          input_mem_banks_bank_a_35_sva_dfm_2, input_mem_banks_bank_a_36_sva_dfm_2,
          input_mem_banks_bank_a_37_sva_dfm_2, input_mem_banks_bank_a_38_sva_dfm_2,
          input_mem_banks_bank_a_39_sva_dfm_2, input_mem_banks_bank_a_40_sva_dfm_2,
          input_mem_banks_bank_a_41_sva_dfm_2, input_mem_banks_bank_a_42_sva_dfm_2,
          input_mem_banks_bank_a_43_sva_dfm_2, input_mem_banks_bank_a_44_sva_dfm_2,
          input_mem_banks_bank_a_45_sva_dfm_2, input_mem_banks_bank_a_46_sva_dfm_2,
          input_mem_banks_bank_a_47_sva_dfm_2, input_mem_banks_bank_a_48_sva_dfm_2,
          input_mem_banks_bank_a_49_sva_dfm_2, input_mem_banks_bank_a_50_sva_dfm_2,
          input_mem_banks_bank_a_51_sva_dfm_2, input_mem_banks_bank_a_52_sva_dfm_2,
          input_mem_banks_bank_a_53_sva_dfm_2, input_mem_banks_bank_a_54_sva_dfm_2,
          input_mem_banks_bank_a_55_sva_dfm_2, input_mem_banks_bank_a_56_sva_dfm_2,
          input_mem_banks_bank_a_57_sva_dfm_2, input_mem_banks_bank_a_58_sva_dfm_2,
          input_mem_banks_bank_a_59_sva_dfm_2, input_mem_banks_bank_a_60_sva_dfm_2,
          input_mem_banks_bank_a_61_sva_dfm_2, input_mem_banks_bank_a_62_sva_dfm_2,
          input_mem_banks_bank_a_63_sva_dfm_2, input_mem_banks_bank_a_64_sva_dfm_2,
          input_mem_banks_bank_a_65_sva_dfm_2, input_mem_banks_bank_a_66_sva_dfm_2,
          input_mem_banks_bank_a_67_sva_dfm_2, input_mem_banks_bank_a_68_sva_dfm_2,
          input_mem_banks_bank_a_69_sva_dfm_2, input_mem_banks_bank_a_70_sva_dfm_2,
          input_mem_banks_bank_a_71_sva_dfm_2, input_mem_banks_bank_a_72_sva_dfm_2,
          input_mem_banks_bank_a_73_sva_dfm_2, input_mem_banks_bank_a_74_sva_dfm_2,
          input_mem_banks_bank_a_75_sva_dfm_2, input_mem_banks_bank_a_76_sva_dfm_2,
          input_mem_banks_bank_a_77_sva_dfm_2, input_mem_banks_bank_a_78_sva_dfm_2,
          input_mem_banks_bank_a_79_sva_dfm_2, input_mem_banks_bank_a_80_sva_dfm_2,
          input_mem_banks_bank_a_81_sva_dfm_2, input_mem_banks_bank_a_82_sva_dfm_2,
          input_mem_banks_bank_a_83_sva_dfm_2, input_mem_banks_bank_a_84_sva_dfm_2,
          input_mem_banks_bank_a_85_sva_dfm_2, input_mem_banks_bank_a_86_sva_dfm_2,
          input_mem_banks_bank_a_87_sva_dfm_2, input_mem_banks_bank_a_88_sva_dfm_2,
          input_mem_banks_bank_a_89_sva_dfm_2, input_mem_banks_bank_a_90_sva_dfm_2,
          input_mem_banks_bank_a_91_sva_dfm_2, input_mem_banks_bank_a_92_sva_dfm_2,
          input_mem_banks_bank_a_93_sva_dfm_2, input_mem_banks_bank_a_94_sva_dfm_2,
          input_mem_banks_bank_a_95_sva_dfm_2, input_mem_banks_bank_a_96_sva_dfm_2,
          input_mem_banks_bank_a_97_sva_dfm_2, input_mem_banks_bank_a_98_sva_dfm_2,
          input_mem_banks_bank_a_99_sva_dfm_2, input_mem_banks_bank_a_100_sva_dfm_2,
          input_mem_banks_bank_a_101_sva_dfm_2, input_mem_banks_bank_a_102_sva_dfm_2,
          input_mem_banks_bank_a_103_sva_dfm_2, input_mem_banks_bank_a_104_sva_dfm_2,
          input_mem_banks_bank_a_105_sva_dfm_2, input_mem_banks_bank_a_106_sva_dfm_2,
          input_mem_banks_bank_a_107_sva_dfm_2, input_mem_banks_bank_a_108_sva_dfm_2,
          input_mem_banks_bank_a_109_sva_dfm_2, input_mem_banks_bank_a_110_sva_dfm_2,
          input_mem_banks_bank_a_111_sva_dfm_2, input_mem_banks_bank_a_112_sva_dfm_2,
          input_mem_banks_bank_a_113_sva_dfm_2, input_mem_banks_bank_a_114_sva_dfm_2,
          input_mem_banks_bank_a_115_sva_dfm_2, input_mem_banks_bank_a_116_sva_dfm_2,
          input_mem_banks_bank_a_117_sva_dfm_2, input_mem_banks_bank_a_118_sva_dfm_2,
          input_mem_banks_bank_a_119_sva_dfm_2, input_mem_banks_bank_a_120_sva_dfm_2,
          input_mem_banks_bank_a_121_sva_dfm_2, input_mem_banks_bank_a_122_sva_dfm_2,
          input_mem_banks_bank_a_123_sva_dfm_2, input_mem_banks_bank_a_124_sva_dfm_2,
          input_mem_banks_bank_a_125_sva_dfm_2, input_mem_banks_bank_a_126_sva_dfm_2,
          input_mem_banks_bank_a_127_sva_dfm_2, input_mem_banks_bank_a_128_sva_dfm_2,
          input_mem_banks_bank_a_129_sva_dfm_2, input_mem_banks_bank_a_130_sva_dfm_2,
          input_mem_banks_bank_a_131_sva_dfm_2, input_mem_banks_bank_a_132_sva_dfm_2,
          input_mem_banks_bank_a_133_sva_dfm_2, input_mem_banks_bank_a_134_sva_dfm_2,
          input_mem_banks_bank_a_135_sva_dfm_2, input_mem_banks_bank_a_136_sva_dfm_2,
          input_mem_banks_bank_a_137_sva_dfm_2, input_mem_banks_bank_a_138_sva_dfm_2,
          input_mem_banks_bank_a_139_sva_dfm_2, input_mem_banks_bank_a_140_sva_dfm_2,
          input_mem_banks_bank_a_141_sva_dfm_2, input_mem_banks_bank_a_142_sva_dfm_2,
          input_mem_banks_bank_a_143_sva_dfm_2, input_mem_banks_bank_a_144_sva_dfm_2,
          input_mem_banks_bank_a_145_sva_dfm_2, input_mem_banks_bank_a_146_sva_dfm_2,
          input_mem_banks_bank_a_147_sva_dfm_2, input_mem_banks_bank_a_148_sva_dfm_2,
          input_mem_banks_bank_a_149_sva_dfm_2, input_mem_banks_bank_a_150_sva_dfm_2,
          input_mem_banks_bank_a_151_sva_dfm_2, input_mem_banks_bank_a_152_sva_dfm_2,
          input_mem_banks_bank_a_153_sva_dfm_2, input_mem_banks_bank_a_154_sva_dfm_2,
          input_mem_banks_bank_a_155_sva_dfm_2, input_mem_banks_bank_a_156_sva_dfm_2,
          input_mem_banks_bank_a_157_sva_dfm_2, input_mem_banks_bank_a_158_sva_dfm_2,
          input_mem_banks_bank_a_159_sva_dfm_2, input_mem_banks_bank_a_160_sva_dfm_2,
          input_mem_banks_bank_a_161_sva_dfm_2, input_mem_banks_bank_a_162_sva_dfm_2,
          input_mem_banks_bank_a_163_sva_dfm_2, input_mem_banks_bank_a_164_sva_dfm_2,
          input_mem_banks_bank_a_165_sva_dfm_2, input_mem_banks_bank_a_166_sva_dfm_2,
          input_mem_banks_bank_a_167_sva_dfm_2, input_mem_banks_bank_a_168_sva_dfm_2,
          input_mem_banks_bank_a_169_sva_dfm_2, input_mem_banks_bank_a_170_sva_dfm_2,
          input_mem_banks_bank_a_171_sva_dfm_2, input_mem_banks_bank_a_172_sva_dfm_2,
          input_mem_banks_bank_a_173_sva_dfm_2, input_mem_banks_bank_a_174_sva_dfm_2,
          input_mem_banks_bank_a_175_sva_dfm_2, input_mem_banks_bank_a_176_sva_dfm_2,
          input_mem_banks_bank_a_177_sva_dfm_2, input_mem_banks_bank_a_178_sva_dfm_2,
          input_mem_banks_bank_a_179_sva_dfm_2, input_mem_banks_bank_a_180_sva_dfm_2,
          input_mem_banks_bank_a_181_sva_dfm_2, input_mem_banks_bank_a_182_sva_dfm_2,
          input_mem_banks_bank_a_183_sva_dfm_2, input_mem_banks_bank_a_184_sva_dfm_2,
          input_mem_banks_bank_a_185_sva_dfm_2, input_mem_banks_bank_a_186_sva_dfm_2,
          input_mem_banks_bank_a_187_sva_dfm_2, input_mem_banks_bank_a_188_sva_dfm_2,
          input_mem_banks_bank_a_189_sva_dfm_2, input_mem_banks_bank_a_190_sva_dfm_2,
          input_mem_banks_bank_a_191_sva_dfm_2, input_mem_banks_bank_a_192_sva_dfm_2,
          input_mem_banks_bank_a_193_sva_dfm_2, input_mem_banks_bank_a_194_sva_dfm_2,
          input_mem_banks_bank_a_195_sva_dfm_2, input_mem_banks_bank_a_196_sva_dfm_2,
          input_mem_banks_bank_a_197_sva_dfm_2, input_mem_banks_bank_a_198_sva_dfm_2,
          input_mem_banks_bank_a_199_sva_dfm_2, input_mem_banks_bank_a_200_sva_dfm_2,
          input_mem_banks_bank_a_201_sva_dfm_2, input_mem_banks_bank_a_202_sva_dfm_2,
          input_mem_banks_bank_a_203_sva_dfm_2, input_mem_banks_bank_a_204_sva_dfm_2,
          input_mem_banks_bank_a_205_sva_dfm_2, input_mem_banks_bank_a_206_sva_dfm_2,
          input_mem_banks_bank_a_207_sva_dfm_2, input_mem_banks_bank_a_208_sva_dfm_2,
          input_mem_banks_bank_a_209_sva_dfm_2, input_mem_banks_bank_a_210_sva_dfm_2,
          input_mem_banks_bank_a_211_sva_dfm_2, input_mem_banks_bank_a_212_sva_dfm_2,
          input_mem_banks_bank_a_213_sva_dfm_2, input_mem_banks_bank_a_214_sva_dfm_2,
          input_mem_banks_bank_a_215_sva_dfm_2, input_mem_banks_bank_a_216_sva_dfm_2,
          input_mem_banks_bank_a_217_sva_dfm_2, input_mem_banks_bank_a_218_sva_dfm_2,
          input_mem_banks_bank_a_219_sva_dfm_2, input_mem_banks_bank_a_220_sva_dfm_2,
          input_mem_banks_bank_a_221_sva_dfm_2, input_mem_banks_bank_a_222_sva_dfm_2,
          input_mem_banks_bank_a_223_sva_dfm_2, input_mem_banks_bank_a_224_sva_dfm_2,
          input_mem_banks_bank_a_225_sva_dfm_2, input_mem_banks_bank_a_226_sva_dfm_2,
          input_mem_banks_bank_a_227_sva_dfm_2, input_mem_banks_bank_a_228_sva_dfm_2,
          input_mem_banks_bank_a_229_sva_dfm_2, input_mem_banks_bank_a_230_sva_dfm_2,
          input_mem_banks_bank_a_231_sva_dfm_2, input_mem_banks_bank_a_232_sva_dfm_2,
          input_mem_banks_bank_a_233_sva_dfm_2, input_mem_banks_bank_a_234_sva_dfm_2,
          input_mem_banks_bank_a_235_sva_dfm_2, input_mem_banks_bank_a_236_sva_dfm_2,
          input_mem_banks_bank_a_237_sva_dfm_2, input_mem_banks_bank_a_238_sva_dfm_2,
          input_mem_banks_bank_a_239_sva_dfm_2, input_mem_banks_bank_a_240_sva_dfm_2,
          input_mem_banks_bank_a_241_sva_dfm_2, input_mem_banks_bank_a_242_sva_dfm_2,
          input_mem_banks_bank_a_243_sva_dfm_2, input_mem_banks_bank_a_244_sva_dfm_2,
          input_mem_banks_bank_a_245_sva_dfm_2, input_mem_banks_bank_a_246_sva_dfm_2,
          input_mem_banks_bank_a_247_sva_dfm_2, input_mem_banks_bank_a_248_sva_dfm_2,
          input_mem_banks_bank_a_249_sva_dfm_2, input_mem_banks_bank_a_250_sva_dfm_2,
          input_mem_banks_bank_a_251_sva_dfm_2, input_mem_banks_bank_a_252_sva_dfm_2,
          input_mem_banks_bank_a_253_sva_dfm_2, input_mem_banks_bank_a_254_sva_dfm_2,
          input_mem_banks_bank_a_255_sva_dfm_2, input_mem_banks_read_1_for_mux_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_75_nl & while_stage_0_7 ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_6 <= MUX1HOT_s_1_3_2(PECore_RunMac_PECore_RunMac_if_and_svs_5,
          (weight_port_read_out_data_0_7_sva_dfm_mx0w1[7]), PECore_PushAxiRsp_if_else_mux_23_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_40_tmp , while_and_39_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( input_read_req_valid_and_3_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_15_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= 4'b0000;
      rva_out_reg_data_39_36_sva_dfm_4_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_4_1 <= 7'b0000000;
      rva_out_reg_data_62_56_sva_dfm_4_1 <= 7'b0000000;
      rva_out_reg_data_55_48_sva_dfm_4_1 <= 8'b00000000;
    end
    else if ( and_1442_cse ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= MUX1HOT_v_4_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_3_0,
          rva_out_reg_data_35_32_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[35:32]),
          weight_port_read_out_data_0_4_sva_dfm_mx0w2_3_0, {PECore_PushAxiRsp_if_asn_89
          , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_39_36_sva_dfm_4_1 <= MUX1HOT_v_4_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_3_0,
          rva_out_reg_data_39_36_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:36]),
          weight_port_read_out_data_0_4_sva_dfm_mx0w2_7_4, {PECore_PushAxiRsp_if_asn_89
          , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_46_40_sva_dfm_4_1 <= MUX1HOT_v_7_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_6_0,
          rva_out_reg_data_46_40_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[46:40]),
          (weight_port_read_out_data_0_5_sva_dfm_mx0w1[6:0]), {PECore_PushAxiRsp_if_asn_89
          , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_62_56_sva_dfm_4_1 <= MUX1HOT_v_7_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_6_0,
          rva_out_reg_data_62_56_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[62:56]),
          (weight_port_read_out_data_0_7_sva_dfm_mx0w1[6:0]), {PECore_PushAxiRsp_if_asn_89
          , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_55_48_sva_dfm_4_1 <= MUX1HOT_v_8_4_2(rva_out_reg_data_55_48_sva_dfm_1_5,
          rva_out_reg_data_55_48_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_sva_1,
          {PECore_PushAxiRsp_if_asn_89 , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87
          , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_88_sva_dfm_4_1 <= 8'b00000000;
      rva_out_reg_data_79_72_sva_dfm_4_1 <= 8'b00000000;
      rva_out_reg_data_71_64_sva_dfm_4_1 <= 8'b00000000;
      rva_out_reg_data_127_120_sva_dfm_4_1_7_6 <= 2'b00;
      rva_out_reg_data_127_120_sva_dfm_4_1_5_0 <= 6'b000000;
      rva_out_reg_data_119_112_sva_dfm_4_1_7 <= 1'b0;
      rva_out_reg_data_119_112_sva_dfm_4_1_6_0 <= 7'b0000000;
      rva_out_reg_data_111_104_sva_dfm_4_1_7 <= 1'b0;
      rva_out_reg_data_111_104_sva_dfm_4_1_6_0 <= 7'b0000000;
      rva_out_reg_data_103_96_sva_dfm_4_1_7_4 <= 4'b0000;
      rva_out_reg_data_103_96_sva_dfm_4_1_3_0 <= 4'b0000;
      rva_out_reg_data_87_80_sva_dfm_4_1_7_4 <= 4'b0000;
      rva_out_reg_data_87_80_sva_dfm_4_1_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_78_ssc ) begin
      rva_out_reg_data_95_88_sva_dfm_4_1 <= MUX1HOT_v_8_3_2(rva_out_reg_data_95_88_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000,
          weight_port_read_out_data_6_10_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_79_72_sva_dfm_4_1 <= MUX1HOT_v_8_3_2(rva_out_reg_data_79_72_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
          weight_port_read_out_data_6_8_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_71_64_sva_dfm_4_1 <= MUX1HOT_v_8_3_2(rva_out_reg_data_71_64_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
          weight_port_read_out_data_6_7_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_127_120_sva_dfm_4_1_7_6 <= MUX1HOT_v_2_3_2(rva_out_reg_data_127_120_sva_dfm_4_mx0w0_7_6,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000[7:6]),
          (weight_port_read_out_data_6_6_sva_dfm_1[7:6]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_127_120_sva_dfm_4_1_5_0 <= MUX1HOT_v_6_3_2(rva_out_reg_data_127_120_sva_dfm_4_mx0w0_5_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000[5:0]),
          (weight_port_read_out_data_6_6_sva_dfm_1[5:0]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_119_112_sva_dfm_4_1_7 <= MUX1HOT_s_1_3_2(rva_out_reg_data_119_112_sva_dfm_4_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000[7]),
          (weight_port_read_out_data_6_5_sva_dfm_1[7]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_119_112_sva_dfm_4_1_6_0 <= MUX1HOT_v_7_3_2(rva_out_reg_data_119_112_sva_dfm_4_mx0w0_6_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000[6:0]),
          (weight_port_read_out_data_6_5_sva_dfm_1[6:0]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_111_104_sva_dfm_4_1_7 <= MUX1HOT_s_1_3_2(rva_out_reg_data_111_104_sva_dfm_4_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000[7]),
          (weight_port_read_out_data_6_4_sva_dfm_1[7]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_111_104_sva_dfm_4_1_6_0 <= MUX1HOT_v_7_3_2(rva_out_reg_data_111_104_sva_dfm_4_mx0w0_6_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000[6:0]),
          (weight_port_read_out_data_6_4_sva_dfm_1[6:0]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_103_96_sva_dfm_4_1_7_4 <= MUX1HOT_v_4_3_2((rva_out_reg_data_103_96_sva_dfm_4_mx0w0[7:4]),
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005[7:4]),
          weight_port_read_out_data_0_10_sva_dfm_2_7_4, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1243_cse , while_while_nor_259_cse});
      rva_out_reg_data_103_96_sva_dfm_4_1_3_0 <= MUX1HOT_v_4_3_2((rva_out_reg_data_103_96_sva_dfm_4_mx0w0[3:0]),
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005[3:0]),
          weight_port_read_out_data_0_10_sva_dfm_2_3_0, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1243_cse , while_while_nor_259_cse});
      rva_out_reg_data_87_80_sva_dfm_4_1_7_4 <= MUX1HOT_v_4_3_2(rva_out_reg_data_87_80_sva_dfm_4_mx0w0_7_4,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[7:4]),
          (weight_port_read_out_data_6_9_sva_dfm_1[7:4]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
      rva_out_reg_data_87_80_sva_dfm_4_1_3_0 <= MUX1HOT_v_4_3_2(rva_out_reg_data_87_80_sva_dfm_4_mx0w0_3_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[3:0]),
          (weight_port_read_out_data_6_9_sva_dfm_1[3:0]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_552 , and_dcpl_553});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & or_tmp_85 & and_dcpl_40 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_63_sva_dfm_6 <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse & (~ mux_81_nl) ) begin
      rva_out_reg_data_63_sva_dfm_6 <= rva_out_reg_data_63_sva_dfm_6_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_62_56_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_46_40_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_39_36_sva_dfm_6 <= 4'b0000;
      rva_out_reg_data_35_32_sva_dfm_6 <= 4'b0000;
    end
    else if ( and_1463_cse ) begin
      rva_out_reg_data_55_48_sva_dfm_6 <= rva_out_reg_data_55_48_sva_dfm_6_mx1;
      rva_out_reg_data_62_56_sva_dfm_6 <= rva_out_reg_data_62_56_sva_dfm_6_mx1;
      rva_out_reg_data_46_40_sva_dfm_6 <= rva_out_reg_data_46_40_sva_dfm_6_mx1;
      rva_out_reg_data_39_36_sva_dfm_6 <= rva_out_reg_data_39_36_sva_dfm_6_mx1;
      rva_out_reg_data_35_32_sva_dfm_6 <= rva_out_reg_data_35_32_sva_dfm_6_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(rva_in_reg_rw_sva_5 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        | (~ while_stage_0_7))) ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          (weight_port_read_out_data_0_5_sva_dfm_mx0w1[7]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~((~((~ rva_in_reg_rw_sva_st_1_4) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1
        & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2))) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
        & while_stage_0_6 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= MUX1HOT_v_128_3_2(input_mem_banks_read_read_data_lpi_1_dfm_1_3,
          weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d, weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1,
          {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          , and_667_nl , nor_499_nl});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_5 <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_82_nl & and_dcpl_54 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_5 <= MUX_v_8_2_2(rva_out_reg_data_55_48_sva_dfm_1_4,
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_79_72_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_95_88_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_103_96_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_111_104_sva_dfm_6_6_0 <= 7'b0000000;
      rva_out_reg_data_119_112_sva_dfm_6_6_0 <= 7'b0000000;
      rva_out_reg_data_127_120_sva_dfm_6_5_0 <= 6'b000000;
      rva_out_reg_data_87_80_sva_dfm_6_7_4 <= 4'b0000;
      rva_out_reg_data_87_80_sva_dfm_6_3_0 <= 4'b0000;
    end
    else if ( and_1488_cse ) begin
      rva_out_reg_data_71_64_sva_dfm_6 <= rva_out_reg_data_71_64_sva_dfm_4_mx0w0;
      rva_out_reg_data_79_72_sva_dfm_6 <= rva_out_reg_data_79_72_sva_dfm_4_mx0w0;
      rva_out_reg_data_95_88_sva_dfm_6 <= rva_out_reg_data_95_88_sva_dfm_4_mx0w0;
      rva_out_reg_data_103_96_sva_dfm_6 <= rva_out_reg_data_103_96_sva_dfm_4_mx0w0;
      rva_out_reg_data_111_104_sva_dfm_6_6_0 <= rva_out_reg_data_111_104_sva_dfm_4_mx0w0_6_0;
      rva_out_reg_data_119_112_sva_dfm_6_6_0 <= rva_out_reg_data_119_112_sva_dfm_4_mx0w0_6_0;
      rva_out_reg_data_127_120_sva_dfm_6_5_0 <= rva_out_reg_data_127_120_sva_dfm_4_mx0w0_5_0;
      rva_out_reg_data_87_80_sva_dfm_6_7_4 <= rva_out_reg_data_87_80_sva_dfm_4_mx0w0_7_4;
      rva_out_reg_data_87_80_sva_dfm_6_3_0 <= rva_out_reg_data_87_80_sva_dfm_4_mx0w0_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_221_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_221_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_225_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_225_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_229_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_229_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_233_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_233_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_237_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_237_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_241_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_241_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_245_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_245_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_249_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_249_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_253_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_253_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_257_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_257_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_261_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_261_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_265_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_265_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_269_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_269_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_273_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_273_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_277_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_277_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_281_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_281_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_285_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_285_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_289_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_289_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_293_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_293_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_297_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_297_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_301_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_301_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_305_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_305_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_309_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_309_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_313_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_313_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_317_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_317_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_321_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_321_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_325_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_325_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_329_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_329_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_333_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_333_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_337_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_337_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_341_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_341_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_345_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_345_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_349_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_349_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_353_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_353_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_357_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_357_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_361_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_361_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_365_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_365_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_369_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_369_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_373_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_373_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_377_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_377_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_381_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_381_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_385_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_385_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_389_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_389_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_393_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_393_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_397_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_397_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_401_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_401_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_405_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_405_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_409_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_409_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_413_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_413_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_417_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_417_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_421_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_421_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_425_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_425_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_429_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_429_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_433_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_433_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_437_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_437_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_441_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_441_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_445_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_445_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_449_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_449_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_453_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_453_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_457_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_457_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_461_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_461_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_465_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_465_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_469_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_469_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_473_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_473_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_477_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_477_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_481_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_481_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_485_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_485_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_489_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_489_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_493_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_493_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_497_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_497_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_501_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_501_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_505_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_505_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_509_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_509_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_513_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_513_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_517_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_517_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_521_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_521_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_525_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_525_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_529_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_529_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_533_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_533_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_537_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_537_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_541_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_541_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_545_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_545_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_549_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_549_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_553_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_553_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_557_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_557_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_561_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_561_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_565_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_565_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_569_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_569_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_573_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_573_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_577_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_577_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_581_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_581_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_585_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_585_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_589_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_589_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_593_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_593_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_597_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_597_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_601_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_601_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_605_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_605_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_609_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_609_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_613_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_613_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_617_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_617_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_621_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_621_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_625_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_625_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_629_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_629_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_633_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_633_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_637_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_637_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_641_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_641_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_645_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_645_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_649_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_649_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_653_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_653_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_657_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_657_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_661_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_661_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_665_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_665_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_669_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_669_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_673_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_673_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_677_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_677_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_681_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_681_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_685_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_685_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_689_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_689_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_693_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_693_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_697_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_697_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_701_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_701_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_705_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_705_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_709_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_709_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_713_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_713_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_717_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_717_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_721_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_721_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_725_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_725_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_729_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_729_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_733_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_733_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_737_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_737_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_741_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_741_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_745_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_745_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_749_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_749_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_753_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_753_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_757_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_757_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_761_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_761_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_765_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_765_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_769_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_769_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_773_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_773_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_777_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_777_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_781_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_781_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_785_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_785_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_789_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_789_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_793_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_793_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_797_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_797_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_801_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_801_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_805_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_805_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_809_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_809_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_813_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_813_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_817_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_817_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_821_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_821_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_825_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_825_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_829_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_829_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_833_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_833_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_837_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_837_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_841_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_841_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_845_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_845_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_849_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_849_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_853_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_853_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_857_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_857_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_861_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_861_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_865_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_865_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_869_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_869_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_873_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_873_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_877_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_877_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_881_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_881_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_885_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_885_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_889_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_889_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_893_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_893_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_897_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_897_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_901_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_901_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_905_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_905_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_909_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_909_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_913_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_913_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_917_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_917_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_921_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_921_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_925_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_925_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_929_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_929_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_933_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_933_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_937_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_937_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_941_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_941_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_945_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_945_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_949_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_949_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_953_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_953_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_957_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_957_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_961_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_961_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_965_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_965_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_969_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_969_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_973_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_973_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_977_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_977_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_981_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_981_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_985_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_985_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_989_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_989_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_993_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_993_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_997_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_997_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1001_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1001_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1005_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1005_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1009_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1009_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1013_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1013_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1017_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1017_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1021_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1021_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1025_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1025_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1029_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1029_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1033_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1033_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1037_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1037_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1041_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1041_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1045_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1045_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1049_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1049_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1053_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1053_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1057_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1057_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1061_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1061_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1065_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1065_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1069_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1069_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1073_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1073_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1077_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1077_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1081_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1081_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1085_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1085_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1089_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1089_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1093_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1093_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1097_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1097_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1101_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1101_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1105_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1105_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1109_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1109_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1113_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1113_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1117_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1117_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1121_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1121_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1125_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1125_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1129_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1129_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1133_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1133_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1137_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1137_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1141_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1141_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1145_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1145_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1149_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1149_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1153_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1153_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1157_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1157_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1161_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1161_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1165_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1165_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1169_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1169_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1173_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1173_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1177_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1177_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1181_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1181_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1185_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1185_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1189_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1189_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1193_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1193_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1197_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1197_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1201_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1201_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1205_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1205_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1209_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1209_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1213_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1213_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1217_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1217_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1221_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1221_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1225_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1225_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1229_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1229_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1233_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1233_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1237_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1237_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1241_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1241_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_91_nl) & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_5 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_10_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_5 <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_19_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_base_input_and_tmp ) begin
      pe_manager_base_input_sva <= MUX_v_15_2_2(pe_manager_base_input_sva_dfm_3_1,
          while_if_while_if_and_2_nl, and_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_sva_1_load <= 1'b1;
      accum_vector_data_6_sva_1_load <= 1'b1;
      accum_vector_data_5_sva_1_load <= 1'b1;
      accum_vector_data_3_sva_1_load <= 1'b1;
      accum_vector_data_1_sva_1_load <= 1'b1;
      accum_vector_data_0_sva_1_load <= 1'b1;
      accum_vector_data_4_sva_1_load <= 1'b1;
      accum_vector_data_2_sva_1_load <= 1'b1;
    end
    else if ( and_724_cse ) begin
      accum_vector_data_7_sva_1_load <= accum_vector_data_7_sva_1_load_mx0w1 & (~
          and_dcpl_663);
      accum_vector_data_6_sva_1_load <= accum_vector_data_6_sva_1_load_mx0w1 & (~
          and_dcpl_663);
      accum_vector_data_5_sva_1_load <= accum_vector_data_5_sva_1_load_mx0w0 & (~
          and_dcpl_663);
      accum_vector_data_3_sva_1_load <= accum_vector_data_3_sva_1_load_mx0w1 & (~
          and_dcpl_663);
      accum_vector_data_1_sva_1_load <= accum_vector_data_1_sva_1_load_mx0w1 & (~
          and_dcpl_663);
      accum_vector_data_0_sva_1_load <= accum_vector_data_0_sva_1_load_mx0w1 & (~
          and_dcpl_663);
      accum_vector_data_4_sva_1_load <= accum_vector_data_4_sva_1_load_mx0w0 & (~
          and_dcpl_663);
      accum_vector_data_2_sva_1_load <= accum_vector_data_2_sva_1_load_mx0w0 & (~
          and_dcpl_663);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( (~((~((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6:4]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:7]!=3'b000))) & nor_589_cse
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:12]!=3'b000))) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]))
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & rva_in_PopNB_mioi_return_rsc_z_mxwt
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]==2'b00) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt))
        & while_stage_0_3)) & rva_in_reg_rw_and_5_cse ) begin
      pe_manager_base_input_sva_dfm_3_1 <= MUX_v_15_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[62:48]),
          pe_manager_base_input_sva_mx2, or_512_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & ((nor_384_cse & while_stage_0_3) | and_dcpl_497) )
        begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_operator_1_for_asn_73_itm_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(reg_rva_in_reg_rw_sva_2_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      accum_vector_operator_1_for_asn_73_itm_2 <= accum_vector_operator_1_for_asn_73_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_operator_1_for_asn_43_itm_2 <= 1'b0;
      accum_vector_operator_1_for_asn_28_itm_2 <= 1'b0;
    end
    else if ( accum_vector_operator_1_for_and_45_cse ) begin
      accum_vector_operator_1_for_asn_43_itm_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
      accum_vector_operator_1_for_asn_28_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_94_nl & while_stage_0_5 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= MUX_s_1_2_2((pe_manager_base_weight_sva[0]), PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_3 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_33_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_23_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          accum_vector_operator_1_for_asn_28_itm_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          accum_vector_operator_1_for_asn_43_itm_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_168_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= rva_out_reg_data_30_25_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_169_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= rva_out_reg_data_23_17_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_170_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= rva_out_reg_data_15_9_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_171_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= rva_out_reg_data_35_32_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_172_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= rva_out_reg_data_39_36_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_173_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= rva_out_reg_data_46_40_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_174_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_4 <= rva_out_reg_data_62_56_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_175_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_4 <= rva_out_reg_data_55_48_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]))) & while_stage_0_4 )
        begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_operator_1_for_asn_73_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        & while_stage_0_3 ) begin
      accum_vector_operator_1_for_asn_73_itm_1 <= MUX_s_1_2_2(accum_vector_data_4_sva_1_load_mx0w0,
          ProductSum_for_asn_56_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_96_nl) & while_stage_0_4 ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_3 <= MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_34_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= 6'b000000;
      rva_out_reg_data_23_17_sva_dfm_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_109_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= MUX_v_6_2_2(6'b000000, (pe_manager_base_weight_sva_mx2[14:9]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
      rva_out_reg_data_23_17_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_base_weight_sva_mx2[7:1]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_176_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= rva_out_reg_data_15_9_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_177_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= rva_out_reg_data_35_32_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_178_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= rva_out_reg_data_39_36_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_179_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= rva_out_reg_data_46_40_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_180_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_3 <= rva_out_reg_data_62_56_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_181_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_3 <= rva_out_reg_data_55_48_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_97_nl) & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_29_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= MUX_s_1_2_2(accum_vector_data_1_sva_1_load_mx0w1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_2_1,
          PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= MUX_s_1_2_2(accum_vector_data_2_sva_1_load_mx0w0,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_117_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= rva_out_reg_data_15_9_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_182_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= rva_out_reg_data_35_32_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_183_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= rva_out_reg_data_39_36_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_184_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= rva_out_reg_data_46_40_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_185_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_2 <= rva_out_reg_data_62_56_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_186_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_2 <= pe_config_input_counter_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~(and_dcpl_477 & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[2])
        & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_1 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2))
        & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3) & PECore_DecodeAxiRead_switch_lp_nor_2_cse))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        & while_stage_0_3 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= MUX_s_1_2_2(accum_vector_data_7_sva_1_load_mx0w1,
          PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= MUX_s_1_2_2(accum_vector_data_0_sva_1_load_mx0w1,
          PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(accum_vector_data_6_sva_1_load_mx0w1,
          PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_35_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_497 ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_2 <= PECore_RunMac_PECore_RunMac_if_and_svs_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_1 <= 7'b0000000;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0);
      rva_out_reg_data_15_9_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_num_input_sva[7:1]),
          and_315_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_40_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= pe_config_is_cluster_sva;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1 <= pe_config_is_bias_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= 1'b0;
      rva_out_reg_data_35_32_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_39_36_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_1_1 <= 7'b0000000;
      rva_out_reg_data_62_56_sva_dfm_1_1 <= 7'b0000000;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= (pe_config_num_output_sva[7]) & (~(and_315_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0))
          & PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
      rva_out_reg_data_35_32_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl
          & (signext_4_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0))
          & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_39_36_sva_dfm_1_1 <= (pe_manager_base_bias_sva[7:4]) & ({{3{and_315_cse}},
          and_315_cse}) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_46_40_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl
          & (signext_7_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0))
          & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_62_56_sva_dfm_1_1 <= (pe_manager_base_input_sva_mx2[14:8])
          & ({{6{and_315_cse}}, and_315_cse}) & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_5_mux_107_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_107_itm_1_6_0 <= 7'b0000000;
      weight_mem_run_3_for_5_mux_109_itm_1_7_6 <= 2'b00;
      weight_mem_run_3_for_5_mux_109_itm_1_5_0 <= 6'b000000;
      weight_mem_run_3_for_5_mux_108_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_108_itm_1_6_0 <= 7'b0000000;
      weight_mem_run_3_for_5_mux_11_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_11_itm_1_6_0 <= 7'b0000000;
    end
    else if ( weight_mem_run_3_for_5_and_199_ssc ) begin
      weight_mem_run_3_for_5_mux_107_itm_1_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[7]),
          (weight_port_read_out_data_6_11_sva_dfm_1[7]), and_dcpl_553);
      weight_mem_run_3_for_5_mux_107_itm_1_6_0 <= MUX1HOT_v_7_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[6:0]),
          (weight_port_read_out_data_6_11_sva_dfm_1[6:0]), (input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:9]),
          {and_dcpl_552 , and_dcpl_553 , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
      weight_mem_run_3_for_5_mux_109_itm_1_7_6 <= MUX_v_2_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[7:6]),
          (weight_port_read_out_data_6_13_sva_dfm_1[7:6]), and_dcpl_553);
      weight_mem_run_3_for_5_mux_109_itm_1_5_0 <= MUX1HOT_v_6_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[5:0]),
          (weight_port_read_out_data_6_13_sva_dfm_1[5:0]), (input_mem_banks_read_read_data_lpi_1_dfm_1_4[30:25]),
          {and_dcpl_552 , and_dcpl_553 , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
      weight_mem_run_3_for_5_mux_108_itm_1_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[7]),
          (weight_port_read_out_data_6_12_sva_dfm_1[7]), and_dcpl_553);
      weight_mem_run_3_for_5_mux_108_itm_1_6_0 <= MUX1HOT_v_7_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[6:0]),
          (weight_port_read_out_data_6_12_sva_dfm_1[6:0]), (input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:17]),
          {and_dcpl_552 , and_dcpl_553 , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
      weight_mem_run_3_for_5_mux_11_itm_1_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004[7]),
          (weight_port_read_out_data_0_11_sva_dfm_2[7]), while_while_nor_259_cse);
      weight_mem_run_3_for_5_mux_11_itm_1_6_0 <= MUX1HOT_v_7_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004[6:0]),
          (weight_port_read_out_data_0_11_sva_dfm_2[6:0]), (input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:1]),
          {while_and_1243_cse , while_while_nor_259_cse , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_5_mux_111_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_111_itm_1_6_0 <= 7'b0000000;
      weight_mem_run_3_for_5_mux_110_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_110_itm_1_6_0 <= 7'b0000000;
      weight_mem_run_3_for_5_mux_12_itm_1_7_6 <= 2'b00;
      weight_mem_run_3_for_5_mux_12_itm_1_5_0 <= 6'b000000;
    end
    else if ( weight_mem_run_3_for_5_and_202_ssc ) begin
      weight_mem_run_3_for_5_mux_111_itm_1_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[7]),
          (weight_port_read_out_data_6_15_sva_dfm_1[7]), and_dcpl_553);
      weight_mem_run_3_for_5_mux_111_itm_1_6_0 <= MUX1HOT_v_7_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[6:0]),
          (weight_port_read_out_data_6_15_sva_dfm_1[6:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0,
          {and_dcpl_552 , and_dcpl_553 , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
      weight_mem_run_3_for_5_mux_110_itm_1_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[7]),
          (weight_port_read_out_data_6_14_sva_dfm_1[7]), and_dcpl_553);
      weight_mem_run_3_for_5_mux_110_itm_1_6_0 <= MUX1HOT_v_7_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000[6:0]),
          (weight_port_read_out_data_6_14_sva_dfm_1[6:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0,
          {and_dcpl_552 , and_dcpl_553 , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
      weight_mem_run_3_for_5_mux_12_itm_1_7_6 <= MUX_v_2_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007[7:6]),
          (weight_port_read_out_data_0_12_sva_dfm_2[7:6]), while_while_nor_259_cse);
      weight_mem_run_3_for_5_mux_12_itm_1_5_0 <= MUX1HOT_v_6_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007[5:0]),
          (weight_port_read_out_data_0_12_sva_dfm_2[5:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_5_0,
          {while_and_1243_cse , while_while_nor_259_cse , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_7_4 <= 4'b0000;
      weight_port_read_out_data_0_1_sva_dfm_1_3_0 <= 4'b0000;
      weight_port_read_out_data_0_3_sva_dfm_1_6_0 <= 7'b0000000;
    end
    else if ( and_1529_cse ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_7_4 <= MUX_v_4_2_2(4'b0000, mux1h_3_nl,
          not_2368_nl);
      weight_port_read_out_data_0_1_sva_dfm_1_3_0 <= MUX_v_4_2_2(4'b0000, mux1h_15_nl,
          not_2277_nl);
      weight_port_read_out_data_0_3_sva_dfm_1_6_0 <= MUX_v_7_2_2(7'b0000000, mux1h_13_nl,
          not_2366_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_7 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_1_7 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_136_ssc ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_7 <= mux1h_4_nl & (~ or_dcpl);
      weight_port_read_out_data_0_2_sva_dfm_1_7 <= mux1h_5_nl & (~ or_dcpl_329);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_6_0 <= 7'b0000000;
    end
    else if ( and_1538_tmp ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_6_0 <= MUX_v_7_2_2(7'b0000000, mux1h_14_nl,
          not_2367_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_7_4
          <= 4'b0000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_3_0
          <= 4'b0000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_6_0
          <= 7'b0000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_7_4
          <= MUX_v_4_2_2(4'b0000, weight_mem_banks_load_store_for_else_mux1h_3_nl,
          not_2269_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_3_0
          <= MUX_v_4_2_2(4'b0000, weight_mem_banks_load_store_for_else_mux1h_87_nl,
          not_2270_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_76_nl & (~ or_dcpl_331);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_88_nl,
          not_2272_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_81_nl & (~ or_dcpl_331);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_89_nl,
          not_2274_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7_6
          <= 2'b00;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_5_0
          <= 6'b000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0
          <= 7'b0000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_3_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7_6
          <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm[7:6];
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_5_0
          <= MUX_v_6_2_2(rva_out_reg_data_30_25_sva_dfm_2, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm[5:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7
          <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm[7];
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0
          <= MUX_v_7_2_2(rva_out_reg_data_23_17_sva_dfm_2, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm[6:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7
          <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm[7];
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0
          <= MUX_v_7_2_2(rva_out_reg_data_15_9_sva_dfm_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm[6:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7_4
          <= 4'b0000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_3_0
          <= 4'b0000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_77_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7_4
          <= MUX_v_4_2_2(4'b0000, mux_415_nl, not_2275_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_3_0
          <= MUX_v_4_2_2(4'b0000, mux_416_nl, not_2276_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_248_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_0 <= weight_port_read_out_data_0_1_sva_dfm_1_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_249_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_1 <= weight_port_read_out_data_0_1_sva_dfm_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_2_rsp_0 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_209_ssc ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_0 <= weight_port_read_out_data_0_2_sva_dfm_1_7;
      weight_port_read_out_data_0_3_sva_dfm_2_rsp_0 <= weight_port_read_out_data_0_3_sva_dfm_1_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_250_enex5 ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_1 <= weight_port_read_out_data_0_2_sva_dfm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_rsp_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_251_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_rsp_1 <= weight_port_read_out_data_0_3_sva_dfm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_6_3 <=
          4'b0000;
    end
    else if ( weight_port_read_out_data_and_252_enex5 ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_6_3 <=
          reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_5_0 <=
          6'b000000;
    end
    else if ( weight_port_read_out_data_and_253_enex5 ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_5_0 <=
          reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_1[6:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_4_6_0 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_254_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_4_6_0 <= reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_1_7_4 <= 4'b0000;
      weight_port_read_out_data_0_0_sva_dfm_1_1_3_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_129_ssc ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_1_7_4 <= MUX_v_4_2_2(weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_7_4,
          weight_port_read_out_data_0_0_sva_dfm_mx0w1_7_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
      weight_port_read_out_data_0_0_sva_dfm_1_1_3_0 <= MUX_v_4_2_2(weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_3_0,
          weight_port_read_out_data_0_0_sva_dfm_mx0w1_3_0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1_7 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_1_1_7 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_130_ssc ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1_7 <= MUX1HOT_s_1_9_2(weight_port_read_out_data_0_3_sva_mx0_7,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[31]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_cse
          , weight_mem_run_3_for_5_and_157_ssc , weight_mem_run_3_for_5_and_158_ssc
          , weight_mem_run_3_for_5_and_159_cse , weight_mem_run_3_for_5_and_160_ssc
          , weight_mem_run_3_for_5_and_161_cse , weight_mem_run_3_for_5_and_162_ssc
          , weight_mem_run_3_for_5_and_163_ssc});
      weight_port_read_out_data_0_2_sva_dfm_1_1_7 <= MUX1HOT_s_1_9_2(weight_port_read_out_data_0_2_sva_mx0_7,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[23]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_cse
          , weight_mem_run_3_for_5_and_165_ssc , weight_mem_run_3_for_5_and_166_ssc
          , weight_mem_run_3_for_5_and_159_cse , weight_mem_run_3_for_5_and_168_ssc
          , weight_mem_run_3_for_5_and_161_cse , weight_mem_run_3_for_5_and_170_ssc
          , weight_mem_run_3_for_5_and_171_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1_6_0 <= 7'b0000000;
    end
    else if ( mux_545_nl & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1_6_0 <= MUX1HOT_v_7_9_2(weight_port_read_out_data_0_3_sva_mx0_6_0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[30:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[30:24]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[30:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[30:24]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[30:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[30:24]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[30:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[22:16]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_cse
          , weight_mem_run_3_for_5_and_157_ssc , weight_mem_run_3_for_5_and_158_ssc
          , weight_mem_run_3_for_5_and_159_cse , weight_mem_run_3_for_5_and_160_ssc
          , weight_mem_run_3_for_5_and_161_cse , weight_mem_run_3_for_5_and_162_ssc
          , weight_mem_run_3_for_5_and_163_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_6_0 <= 7'b0000000;
    end
    else if ( mux_547_nl & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_6_0 <= MUX1HOT_v_7_9_2(weight_port_read_out_data_0_2_sva_mx0_6_0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[22:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[22:16]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[22:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[22:16]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[22:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[22:16]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[22:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[14:8]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_cse
          , weight_mem_run_3_for_5_and_165_ssc , weight_mem_run_3_for_5_and_166_ssc
          , weight_mem_run_3_for_5_and_159_cse , weight_mem_run_3_for_5_and_168_ssc
          , weight_mem_run_3_for_5_and_161_cse , weight_mem_run_3_for_5_and_170_ssc
          , weight_mem_run_3_for_5_and_171_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_1_7_4 <= 4'b0000;
      weight_port_read_out_data_0_1_sva_dfm_1_1_3_0 <= 4'b0000;
    end
    else if ( and_1551_cse ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_1_7_4 <= MUX1HOT_v_4_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000[7:4]),
          weight_port_read_out_data_0_1_sva_mx0_7_4, weight_port_read_out_data_0_4_sva_dfm_mx0w2_7_4,
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_nl,
          {and_568_ssc , and_569_ssc , and_570_ssc , and_572_cse});
      weight_port_read_out_data_0_1_sva_dfm_1_1_3_0 <= MUX1HOT_v_4_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000[3:0]),
          weight_port_read_out_data_0_1_sva_mx0_3_0, weight_port_read_out_data_0_4_sva_dfm_mx0w2_3_0,
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_134_nl,
          {and_568_ssc , and_569_ssc , and_570_ssc , and_572_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_255_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_0_sva_dfm_2_7_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_256_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1 <= weight_port_read_out_data_0_0_sva_dfm_2_3_0_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7_4 <= 4'b0000;
      weight_port_read_out_data_0_0_sva_dfm_2_3_0 <= 4'b0000;
    end
    else if ( and_1557_cse ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7_4 <= MUX_v_4_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w1_7_4,
          weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_7_4, and_dcpl_40);
      weight_port_read_out_data_0_0_sva_dfm_2_3_0 <= MUX_v_4_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w1_3_0,
          weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_3_0, and_dcpl_40);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7_4_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_257_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7_4_1 <= weight_port_read_out_data_0_0_sva_dfm_1_1_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_3_0_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_258_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_3_0_1 <= weight_port_read_out_data_0_0_sva_dfm_1_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_120_sva_dfm_4_2_rsp_1 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_187_enex5 ) begin
      rva_out_reg_data_127_120_sva_dfm_4_2_rsp_1 <= rva_out_reg_data_127_120_sva_dfm_4_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_119_112_sva_dfm_4_2_rsp_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_188_enex5 ) begin
      rva_out_reg_data_119_112_sva_dfm_4_2_rsp_1 <= rva_out_reg_data_119_112_sva_dfm_4_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_104_sva_dfm_4_2_rsp_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_189_enex5 ) begin
      rva_out_reg_data_111_104_sva_dfm_4_2_rsp_1 <= rva_out_reg_data_111_104_sva_dfm_4_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_104_sva_dfm_6_7 <= 1'b0;
      rva_out_reg_data_119_112_sva_dfm_6_7 <= 1'b0;
      rva_out_reg_data_127_120_sva_dfm_6_7_6 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_93_cse ) begin
      rva_out_reg_data_111_104_sva_dfm_6_7 <= MUX_s_1_2_2(rva_out_reg_data_111_104_sva_dfm_4_mx0w0_7,
          rva_out_reg_data_111_104_sva_dfm_7_7, while_asn_998);
      rva_out_reg_data_119_112_sva_dfm_6_7 <= MUX_s_1_2_2(rva_out_reg_data_119_112_sva_dfm_4_mx0w0_7,
          rva_out_reg_data_119_112_sva_dfm_7_7, while_asn_998);
      rva_out_reg_data_127_120_sva_dfm_6_7_6 <= MUX_v_2_2_2(rva_out_reg_data_127_120_sva_dfm_4_mx0w0_7_6,
          rva_out_reg_data_127_120_sva_dfm_7_7_6, while_asn_998);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_120_sva_dfm_4_4_5_0 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_190_enex5 ) begin
      rva_out_reg_data_127_120_sva_dfm_4_4_5_0 <= reg_rva_out_reg_data_127_120_sva_dfm_4_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_119_112_sva_dfm_4_4_6_0 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_191_enex5 ) begin
      rva_out_reg_data_119_112_sva_dfm_4_4_6_0 <= reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_104_sva_dfm_4_4_6_0 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_192_enex5 ) begin
      rva_out_reg_data_111_104_sva_dfm_4_4_6_0 <= reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_4_sva_dfm_1_1_7_4 <= 4'b0000;
      weight_port_read_out_data_0_4_sva_dfm_1_1_3_0 <= 4'b0000;
    end
    else if ( and_1580_cse ) begin
      weight_port_read_out_data_0_4_sva_dfm_1_1_7_4 <= MUX1HOT_v_4_9_2(weight_port_read_out_data_0_4_sva_mx0_7_4,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:36]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:36]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:36]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:36]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:36]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:36]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:36]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:28]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_cse
          , weight_mem_run_3_for_5_and_173_cse , weight_mem_run_3_for_5_and_174_cse
          , weight_mem_run_3_for_5_and_159_cse , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_161_cse , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_187_ssc});
      weight_port_read_out_data_0_4_sva_dfm_1_1_3_0 <= MUX1HOT_v_4_9_2(weight_port_read_out_data_0_4_sva_mx0_3_0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[35:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[35:32]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[35:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[35:32]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[35:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[35:32]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[35:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[27:24]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_cse
          , weight_mem_run_3_for_5_and_173_cse , weight_mem_run_3_for_5_and_174_cse
          , weight_mem_run_3_for_5_and_159_cse , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_161_cse , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_187_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_3_rsp_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_193_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_103_96_sva_dfm_4_2_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_3_rsp_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_194_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_103_96_sva_dfm_4_2_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_87_80_sva_dfm_4_3_rsp_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_195_enex5 ) begin
      rva_out_reg_data_87_80_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_87_80_sva_dfm_4_2_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_87_80_sva_dfm_4_3_rsp_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_196_enex5 ) begin
      rva_out_reg_data_87_80_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_87_80_sva_dfm_4_2_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_2_7_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_197_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_2_7_4 <= rva_out_reg_data_103_96_sva_dfm_4_1_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_2_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_198_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_2_3_0 <= rva_out_reg_data_103_96_sva_dfm_4_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_87_80_sva_dfm_4_2_7_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_199_enex5 ) begin
      rva_out_reg_data_87_80_sva_dfm_4_2_7_4 <= rva_out_reg_data_87_80_sva_dfm_4_1_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_87_80_sva_dfm_4_2_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_200_enex5 ) begin
      rva_out_reg_data_87_80_sva_dfm_4_2_3_0 <= rva_out_reg_data_87_80_sva_dfm_4_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_145_enex5 | rva_out_reg_data_and_128_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= rva_out_reg_data_and_145_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_144_enex5 | rva_out_reg_data_and_129_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= rva_out_reg_data_and_144_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_143_enex5 | rva_out_reg_data_and_130_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= rva_out_reg_data_and_143_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_193_enex5 | rva_out_reg_data_and_131_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_3_enexo <= rva_out_reg_data_and_193_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_194_enex5 | rva_out_reg_data_and_132_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_194_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_154_enex5 | rva_out_reg_data_and_133_enex5 ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_enexo <= rva_out_reg_data_and_154_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_195_enex5 | rva_out_reg_data_and_134_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_enexo <= rva_out_reg_data_and_195_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_196_enex5 | rva_out_reg_data_and_135_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_196_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_155_enex5 | rva_out_reg_data_and_136_enex5 ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_3_enexo <= rva_out_reg_data_and_155_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_156_enex5 | rva_out_reg_data_and_137_enex5 ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_3_enexo <= rva_out_reg_data_and_156_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_149_enex5 | rva_out_reg_data_and_138_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo <= rva_out_reg_data_and_149_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_146_enex5 | rva_out_reg_data_and_139_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= rva_out_reg_data_and_146_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_150_enex5 | rva_out_reg_data_and_140_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo <= rva_out_reg_data_and_150_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_147_enex5 | rva_out_reg_data_and_141_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo <= rva_out_reg_data_and_147_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_148_enex5 | rva_out_reg_data_and_142_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo <= rva_out_reg_data_and_148_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_39_enex5 | input_mem_banks_read_read_data_and_35_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo
          <= input_mem_banks_read_read_data_and_39_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_255_enex5 | weight_port_read_out_data_and_213_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_enexo <= weight_port_read_out_data_and_255_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_40_enex5 | input_mem_banks_read_read_data_and_36_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo
          <= input_mem_banks_read_read_data_and_40_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_41_enex5 | input_mem_banks_read_read_data_and_37_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo
          <= input_mem_banks_read_read_data_and_41_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_42_enex5 | input_mem_banks_read_read_data_and_38_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo
          <= input_mem_banks_read_read_data_and_42_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_5_enex5 | input_mem_banks_read_1_read_data_and_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_1_read_data_and_5_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_214_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_215_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_216_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_217_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_218_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_219_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_220_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_221_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_222_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_223_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_224_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_225_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_226_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_227_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_cse | weight_port_read_out_data_and_228_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014
          <= data_in_tmp_operator_2_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_15_tmp | weight_port_read_out_data_and_15_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= data_in_tmp_operator_2_for_and_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_229_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_230_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_231_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_232_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_233_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_234_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_235_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_236_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_237_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_238_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_239_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_240_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_241_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_242_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_243_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_31_tmp | weight_port_read_out_data_and_31_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= data_in_tmp_operator_2_for_and_31_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_6_enex5 | input_mem_banks_read_1_read_data_and_5_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= input_mem_banks_read_1_read_data_and_6_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( weight_read_addrs_and_7_cse | weight_read_addrs_and_28_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= weight_read_addrs_and_7_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_3_lpi_1_dfm_1_enexo <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_weight_read_addrs_3_lpi_1_dfm_1_enexo <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= 1'b1;
    end
    else if ( weight_read_addrs_and_7_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= weight_read_addrs_and_7_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_25_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_3_lpi_1_dfm_1_enexo_1 <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_weight_read_addrs_3_lpi_1_dfm_1_enexo_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= 1'b1;
    end
    else if ( weight_read_addrs_and_7_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= weight_read_addrs_and_7_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= 1'b1;
    end
    else if ( operator_15_false_1_and_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= operator_15_false_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_25_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_64_enex5 | weight_write_data_data_and_48_enex5
        ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_64_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_65_enex5 | weight_write_data_data_and_49_enex5
        ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_65_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_66_enex5 | weight_write_data_data_and_50_enex5
        ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_67_enex5 | weight_write_data_data_and_51_enex5
        ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_68_enex5 | weight_write_data_data_and_52_enex5
        ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_69_enex5 | weight_write_data_data_and_53_enex5
        ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_70_enex5 | weight_write_data_data_and_54_enex5
        ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_70_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_71_enex5 | weight_write_data_data_and_55_enex5
        ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_71_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_72_enex5 | weight_write_data_data_and_56_enex5
        ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_72_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_73_enex5 | weight_write_data_data_and_57_enex5
        ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_73_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_74_enex5 | weight_write_data_data_and_58_enex5
        ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_74_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_75_enex5 | weight_write_data_data_and_59_enex5
        ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_75_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_76_enex5 | weight_write_data_data_and_60_enex5
        ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_76_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_77_enex5 | weight_write_data_data_and_61_enex5
        ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_77_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_78_enex5 | weight_write_data_data_and_62_enex5
        ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_78_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_79_enex5 | weight_write_data_data_and_63_enex5
        ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_79_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_write_addrs_and_2_enex5 | weight_write_addrs_and_enex5 ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= weight_write_addrs_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_64_enex5 ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_65_enex5 ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_66_enex5 ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_67_enex5 ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_68_enex5 ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_69_enex5 ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_70_enex5 ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_71_enex5 ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_72_enex5 ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_73_enex5 ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_74_enex5 ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_75_enex5 ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_76_enex5 ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_77_enex5 ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_78_enex5 ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_79_enex5 ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_input_enexo <= 1'b1;
    end
    else if ( pe_manager_base_input_and_tmp | weight_write_addrs_and_2_enex5 ) begin
      reg_pe_manager_base_input_enexo <= pe_manager_base_input_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_read_addrs_and_29_enex5 ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_config_num_output_enexo <= 1'b1;
    end
    else if ( pe_config_num_manager_and_cse | pe_config_UpdateManagerCounter_if_if_and_enex5
        ) begin
      reg_pe_config_num_output_enexo <= pe_config_num_manager_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_248_enex5 | weight_port_read_out_data_and_244_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_enexo <= weight_port_read_out_data_and_248_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_249_enex5 | weight_port_read_out_data_and_245_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_249_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_250_enex5 | weight_port_read_out_data_and_246_enex5
        ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_250_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_data_sva_1_enexo <= 1'b1;
    end
    else if ( rva_in_reg_data_and_tmp | PEManager_15U_PEManagerWrite_and_enex5 )
        begin
      reg_rva_in_reg_data_sva_1_enexo <= rva_in_reg_data_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_43_enex5 | input_mem_banks_read_read_data_and_39_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= input_mem_banks_read_read_data_and_43_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_44_enex5 | input_mem_banks_read_read_data_and_40_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= input_mem_banks_read_read_data_and_44_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_45_enex5 | input_mem_banks_read_read_data_and_41_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= input_mem_banks_read_read_data_and_45_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_46_enex5 | input_mem_banks_read_read_data_and_42_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= input_mem_banks_read_read_data_and_46_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_7_enex5 | input_mem_banks_read_1_read_data_and_6_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_1_read_data_and_7_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_read_addrs_and_30_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_157_enex5 | rva_out_reg_data_and_143_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= rva_out_reg_data_and_157_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_158_enex5 | rva_out_reg_data_and_144_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= rva_out_reg_data_and_158_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_159_enex5 | rva_out_reg_data_and_145_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= rva_out_reg_data_and_159_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_251_enex5 | weight_port_read_out_data_and_247_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_251_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_160_enex5 | rva_out_reg_data_and_146_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= rva_out_reg_data_and_160_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_161_enex5 | rva_out_reg_data_and_147_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo <= rva_out_reg_data_and_161_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_162_enex5 | rva_out_reg_data_and_148_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo <= rva_out_reg_data_and_162_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_163_enex5 | rva_out_reg_data_and_149_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo <= rva_out_reg_data_and_163_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_164_enex5 | rva_out_reg_data_and_150_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo <= rva_out_reg_data_and_164_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_187_enex5 | rva_out_reg_data_and_151_enex5 ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_187_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_188_enex5 | rva_out_reg_data_and_152_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_188_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_189_enex5 | rva_out_reg_data_and_153_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_189_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_165_enex5 | rva_out_reg_data_and_154_enex5 ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_2_enexo <= rva_out_reg_data_and_165_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_166_enex5 | rva_out_reg_data_and_155_enex5 ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_2_enexo <= rva_out_reg_data_and_166_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_167_enex5 | rva_out_reg_data_and_156_enex5 ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_2_enexo <= rva_out_reg_data_and_167_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_xbar_requests_transpose_and_13_cse | weight_mem_write_arbxbar_xbar_for_empty_and_enex5
        ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= weight_mem_read_arbxbar_xbar_requests_transpose_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_11_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_199_ssc | input_mem_banks_read_read_data_and_43_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_11_itm_1_1_enexo <= weight_mem_run_3_for_5_and_199_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_107_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_199_ssc | input_mem_banks_read_read_data_and_44_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_107_itm_1_1_enexo <= weight_mem_run_3_for_5_and_199_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_108_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_199_ssc | input_mem_banks_read_read_data_and_45_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_108_itm_1_1_enexo <= weight_mem_run_3_for_5_and_199_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_109_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_199_ssc | input_mem_banks_read_read_data_and_46_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_109_itm_1_1_enexo <= weight_mem_run_3_for_5_and_199_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp | input_mem_banks_read_1_read_data_and_7_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= input_mem_banks_read_1_read_data_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_12_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_202_ssc | rva_out_reg_data_and_157_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_12_itm_1_1_enexo <= weight_mem_run_3_for_5_and_202_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_111_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_202_ssc | rva_out_reg_data_and_158_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_111_itm_1_1_enexo <= weight_mem_run_3_for_5_and_202_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_110_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_202_ssc | rva_out_reg_data_and_159_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_110_itm_1_1_enexo <= weight_mem_run_3_for_5_and_202_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1442_cse | rva_out_reg_data_and_160_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= and_1442_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1442_cse | rva_out_reg_data_and_161_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo <= and_1442_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1442_cse | rva_out_reg_data_and_162_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo <= and_1442_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1442_cse | rva_out_reg_data_and_163_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo <= and_1442_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1442_cse | rva_out_reg_data_and_164_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo <= and_1442_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_165_enex5 ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_166_enex5 ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_167_enex5 ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_34_enex5 | input_mem_banks_read_read_data_and_33_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_read_data_and_34_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_109_cse | rva_out_reg_data_and_168_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= rva_out_reg_data_and_109_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_109_cse | rva_out_reg_data_and_169_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= rva_out_reg_data_and_109_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_176_enex5 | rva_out_reg_data_and_170_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= rva_out_reg_data_and_176_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_177_enex5 | rva_out_reg_data_and_171_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= rva_out_reg_data_and_177_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_178_enex5 | rva_out_reg_data_and_172_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= rva_out_reg_data_and_178_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_179_enex5 | rva_out_reg_data_and_173_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= rva_out_reg_data_and_179_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_180_enex5 | rva_out_reg_data_and_174_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo <= rva_out_reg_data_and_180_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_181_enex5 | rva_out_reg_data_and_175_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo <= rva_out_reg_data_and_181_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp | input_mem_banks_read_read_data_and_34_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1 <= input_mem_banks_read_1_read_data_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_117_enex5 | rva_out_reg_data_and_176_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= rva_out_reg_data_and_117_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_182_enex5 | rva_out_reg_data_and_177_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= rva_out_reg_data_and_182_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_183_enex5 | rva_out_reg_data_and_178_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= rva_out_reg_data_and_183_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_184_enex5 | rva_out_reg_data_and_179_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= rva_out_reg_data_and_184_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_185_enex5 | rva_out_reg_data_and_180_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo <= rva_out_reg_data_and_185_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_186_enex5 | rva_out_reg_data_and_181_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo <= rva_out_reg_data_and_186_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse | rva_out_reg_data_and_117_enex5
        ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse | rva_out_reg_data_and_182_enex5
        ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse | rva_out_reg_data_and_183_enex5
        ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse | rva_out_reg_data_and_184_enex5
        ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse | rva_out_reg_data_and_185_enex5
        ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_config_input_counter_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( and_1434_tmp | rva_out_reg_data_and_186_enex5 ) begin
      reg_pe_config_input_counter_sva_dfm_1_enexo <= and_1434_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( and_1529_cse | weight_port_read_out_data_and_248_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_enexo <= and_1529_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1529_cse | weight_port_read_out_data_and_249_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo <= and_1529_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1538_tmp | weight_port_read_out_data_and_250_enex5 ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_1_1_enexo <= and_1538_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1529_cse | weight_port_read_out_data_and_251_enex5 ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_1_enexo <= and_1529_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_244_enex5 | weight_port_read_out_data_and_252_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_enexo <= weight_port_read_out_data_and_244_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_246_enex5 | weight_port_read_out_data_and_253_enex5
        ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_246_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_247_enex5 | weight_port_read_out_data_and_254_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_247_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_257_enex5 | weight_port_read_out_data_and_255_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_enexo <= weight_port_read_out_data_and_257_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_258_enex5 | weight_port_read_out_data_and_256_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_258_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_129_ssc | weight_port_read_out_data_and_257_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo <= weight_port_read_out_data_and_129_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_129_ssc | weight_port_read_out_data_and_258_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_1_enexo <= weight_port_read_out_data_and_129_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_187_enex5 ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_1_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_188_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_1_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_189_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_1_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_151_enex5 | rva_out_reg_data_and_190_enex5 ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_151_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_152_enex5 | rva_out_reg_data_and_191_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_152_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_153_enex5 | rva_out_reg_data_and_192_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_153_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_197_enex5 | rva_out_reg_data_and_193_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_2_enexo <= rva_out_reg_data_and_197_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_198_enex5 | rva_out_reg_data_and_194_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_198_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_199_enex5 | rva_out_reg_data_and_195_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_2_enexo <= rva_out_reg_data_and_199_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_200_enex5 | rva_out_reg_data_and_196_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_200_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_197_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_198_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_1_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_199_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_ssc | rva_out_reg_data_and_200_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_1_1_enexo <= rva_out_reg_data_and_78_ssc;
    end
  end
  assign nl_operator_4_false_acc_nl = pe_config_manager_counter_sva_mx1 + 4'b0001;
  assign operator_4_false_acc_nl = nl_operator_4_false_acc_nl[3:0];
  assign pe_config_UpdateManagerCounter_if_not_7_nl = ~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  assign nl_input_read_addrs_sva_1_1  = pe_config_input_counter_sva_mx1 + pe_manager_base_input_sva_mx1_7_0;
  assign PECore_UpdateFSM_switch_lp_not_23_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_not_24_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_not_25_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_not_26_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_not_27_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_not_28_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_not_29_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_not_19_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign accum_vector_operator_1_for_not_39_nl = ~ accum_vector_operator_1_for_asn_118_itm_6;
  assign accum_vector_operator_1_for_not_38_nl = ~ accum_vector_operator_1_for_asn_103_itm_6;
  assign accum_vector_operator_1_for_not_37_nl = ~ accum_vector_operator_1_for_asn_88_itm_6;
  assign accum_vector_operator_1_for_not_36_nl = ~ accum_vector_operator_1_for_asn_58_itm_6;
  assign accum_vector_operator_1_for_not_35_nl = ~ accum_vector_operator_1_for_asn_28_itm_6;
  assign accum_vector_operator_1_for_not_34_nl = ~ accum_vector_operator_1_for_asn_13_itm_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_1_nl = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign weight_mem_run_3_for_5_and_177_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign and_1270_nl = or_931_cse & mux_tmp_427;
  assign and_1269_nl = or_928_cse & mux_tmp_427;
  assign mux_460_nl = MUX_s_1_2_2(and_1270_nl, and_1269_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_run_3_for_5_and_188_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_191_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign and_1275_nl = or_931_cse & mux_tmp_429;
  assign and_1274_nl = or_928_cse & mux_tmp_429;
  assign mux_462_nl = MUX_s_1_2_2(and_1275_nl, and_1274_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_18_nl = MUX_s_1_2_2(or_tmp_24, and_tmp_1, weight_mem_run_3_for_land_7_lpi_1_dfm_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_136_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_134_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_151_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_28_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign or_52_nl = (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])))
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign or_50_nl = (~(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3)) | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_19_nl = MUX_s_1_2_2(or_50_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3,
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1);
  assign mux_20_nl = MUX_s_1_2_2(or_52_nl, mux_19_nl, while_stage_0_5);
  assign or_48_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_21_nl = MUX_s_1_2_2(mux_20_nl, or_48_nl, while_stage_0_6);
  assign nor_347_nl = ~(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 | (~
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3));
  assign mux_22_nl = MUX_s_1_2_2(nor_347_nl, ProductSum_for_asn_128_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_23_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_3, ProductSum_for_asn_28_itm_3,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign nor_559_nl = ~((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign nor_560_nl = ~((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | (~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1)
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1
      | (~ reg_rva_in_reg_rw_sva_st_1_1_cse));
  assign mux_463_nl = MUX_s_1_2_2(nor_559_nl, nor_560_nl, while_stage_0_3);
  assign mux_464_nl = MUX_s_1_2_2(mux_463_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2,
      while_stage_0_4);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl
      = MUX_v_11_2_2(11'b00000000000, PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl
      = MUX_v_4_2_2(4'b0000, pe_config_manager_counter_sva_mx1, PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign and_638_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & and_dcpl_214 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]));
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl = (state_mux_1_cse!=2'b00)
      | state_0_sva_mx1;
  assign PECore_UpdateFSM_switch_lp_or_nl = PECore_UpdateFSM_switch_lp_equal_tmp_6
      | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  assign PECore_UpdateFSM_switch_lp_mux1h_18_nl = MUX1HOT_v_2_3_2((signext_2_1(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl)),
      2'b01, 2'b10, {PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      , PECore_UpdateFSM_switch_lp_or_nl , PECore_RunScale_PECore_RunScale_if_and_1_svs_1});
  assign PECore_UpdateFSM_switch_lp_nor_8_nl = ~(PECore_PushOutput_PECore_PushOutput_if_and_svs_1
      | PECore_UpdateFSM_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_and_1_nl = MUX_v_2_2_2(2'b00, PECore_UpdateFSM_switch_lp_mux1h_18_nl,
      PECore_UpdateFSM_switch_lp_nor_8_nl);
  assign mux_465_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_3_1, nor_571_cse,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_466_nl = MUX_s_1_2_2(and_1600_cse, nor_571_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nl_operator_8_false_acc_sdt_sva_1  = conv_u2s_8_9(pe_config_num_output_sva)
      + 9'b111111111;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_189_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_199_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_202_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_203_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_219_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_229_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_230_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_232_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign or_196_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_246_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_244_itm_1;
  assign mux_34_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_5_lpi_1_dfm_1, or_196_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_195_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_5_lpi_1_dfm_1;
  assign or_194_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp;
  assign mux_35_nl = MUX_s_1_2_2(mux_34_nl, or_195_nl, or_194_nl);
  assign nor_350_nl = ~((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | rva_in_reg_rw_sva_st_1_4);
  assign nand_39_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & rva_in_reg_rw_sva_st_1_4);
  assign mux_36_nl = MUX_s_1_2_2(nor_350_nl, nand_39_nl, weight_mem_run_3_for_land_6_lpi_1_dfm_1_1);
  assign nor_584_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ or_tmp_541));
  assign mux_489_nl = MUX_s_1_2_2(or_tmp_541, nor_584_nl, while_stage_0_6);
  assign mux_490_nl = MUX_s_1_2_2(mux_489_nl, or_tmp_541, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_48_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[7:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl);
  assign nor_355_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_37_nl = MUX_s_1_2_2(nor_355_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_138_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_80_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[7:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_138_nl);
  assign nor_356_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_208_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1));
  assign mux_38_nl = MUX_s_1_2_2(nor_356_nl, or_208_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_247_itm_1);
  assign or_225_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign mux_40_nl = MUX_s_1_2_2(or_237_cse, or_225_nl, weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp);
  assign nor_359_nl = ~((~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]) |
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]))) | mux_40_nl);
  assign nor_360_nl = ~((~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp)
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign mux_41_nl = MUX_s_1_2_2(nor_359_nl, nor_360_nl, or_222_cse);
  assign nand_2_nl = ~((Arbiter_8U_Roundrobin_pick_1_if_1_and_60_tmp | Arbiter_8U_Roundrobin_pick_1_if_1_and_56_tmp)
      & mux_41_nl);
  assign mux_42_nl = MUX_s_1_2_2(nand_2_nl, or_237_cse, Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp);
  assign or_219_nl = (~ or_dcpl_48) | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign or_217_nl = Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp;
  assign mux_39_nl = MUX_s_1_2_2(or_219_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3,
      or_217_nl);
  assign mux_43_nl = MUX_s_1_2_2(mux_42_nl, mux_39_nl, while_stage_0_5);
  assign mux_57_nl = MUX_s_1_2_2(mux_tmp_49, mux_tmp_43, and_742_cse);
  assign mux_54_nl = MUX_s_1_2_2(mux_tmp_47, mux_tmp_42, and_743_cse);
  assign mux_53_nl = MUX_s_1_2_2(mux_tmp_49, mux_tmp_43, weight_mem_read_arbxbar_arbiters_next_1_3_sva);
  assign mux_55_nl = MUX_s_1_2_2(mux_54_nl, mux_53_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign mux_56_nl = MUX_s_1_2_2(mux_55_nl, mux_47_itm, weight_mem_read_arbxbar_arbiters_next_1_2_sva);
  assign mux_58_nl = MUX_s_1_2_2(mux_57_nl, mux_56_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign mux_48_nl = MUX_s_1_2_2(mux_tmp_43, mux_47_itm, and_744_cse);
  assign mux_49_nl = MUX_s_1_2_2(mux_48_nl, Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp,
      weight_mem_read_arbxbar_arbiters_next_1_6_sva);
  assign mux_59_nl = MUX_s_1_2_2(mux_58_nl, mux_49_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign or_233_nl = (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ mux_59_nl);
  assign or_228_nl = (~ or_dcpl_41) | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign or_226_nl = Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp;
  assign mux_44_nl = MUX_s_1_2_2(or_228_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3,
      or_226_nl);
  assign mux_60_nl = MUX_s_1_2_2(or_233_nl, mux_44_nl, while_stage_0_5);
  assign nand_3_nl = ~((Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_34_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_tmp) & (~((~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]))) | (~ while_stage_0_4)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)));
  assign mux_61_nl = MUX_s_1_2_2(nand_3_nl, or_237_cse, Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp);
  assign or_236_nl = (~(and_745_cse | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp)) |
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_62_nl = MUX_s_1_2_2(mux_61_nl, or_236_nl, while_stage_0_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl
      = pe_manager_base_input_sva_mx1_7_0 & ({{7{and_315_cse}}, and_315_cse}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_1_nl
      = MUX_v_8_2_2(8'b00000000, pe_config_input_counter_sva_mx1, PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl
      = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]), pe_config_is_zero_first_sva_mx1,
      PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_27_nl
      = MUX_s_1_2_2(PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl,
      pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_or_5_cse_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_135_nl = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b101)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_142_nl = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_132_nl = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b110)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b011)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_250_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_175_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_190_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_205_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_220_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_251_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_176_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_191_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_206_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_221_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_252_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_177_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_192_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_207_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_222_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_253_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_178_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_193_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_208_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_223_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_254_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_179_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_194_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_209_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_224_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_255_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_180_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_195_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_210_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_225_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_241_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_181_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_196_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_211_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_226_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_242_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_257_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_182_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_197_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_212_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_227_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_243_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_183_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_198_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_213_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_228_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_238_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[103:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_238_nl);
  assign nor_594_nl = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_2 | (~ and_tmp_17));
  assign mux_495_nl = MUX_s_1_2_2(and_tmp_17, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_496_nl = MUX_s_1_2_2(nor_594_nl, mux_495_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_497_nl = MUX_s_1_2_2(and_tmp_17, mux_496_nl, while_stage_0_6);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_239_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[95:88]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_239_nl);
  assign nor_595_nl = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_2 | (~ and_tmp_18));
  assign mux_501_nl = MUX_s_1_2_2(and_tmp_18, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_502_nl = MUX_s_1_2_2(nor_595_nl, mux_501_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_503_nl = MUX_s_1_2_2(and_tmp_18, mux_502_nl, while_stage_0_6);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_244_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_245_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_247_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_248_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign mux1h_6_nl = MUX1HOT_v_8_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[63:56]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[63:56]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[63:56]),
      {and_1030_cse , and_1031_cse , and_1032_cse});
  assign not_2283_nl = ~ or_dcpl_333;
  assign mux1h_7_nl = MUX1HOT_v_8_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[47:40]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[47:40]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[47:40]),
      {and_1030_cse , and_1031_cse , and_1032_cse});
  assign not_2285_nl = ~ or_dcpl_333;
  assign mux1h_8_nl = MUX1HOT_v_8_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[39:32]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[39:32]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[39:32]),
      {and_1030_cse , and_1031_cse , and_1032_cse});
  assign not_2287_nl = ~ or_dcpl_333;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_200_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_201_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_246_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_140_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_231_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_233_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_port_read_out_data_mux_106_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_23_mx0w2,
      (weight_port_read_out_data_0_7_sva_dfm_mx0w1[7]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1!=3'b000));
  assign mux_73_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, (~ pe_manager_base_weight_slc_pe_manager_base_weight_2_0_371_itm_1),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign nor_371_nl = ~(rva_in_reg_rw_sva_st_1_6 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6));
  assign nor_16_nl = ~(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_6));
  assign mux_74_nl = MUX_s_1_2_2(nand_41_cse, nor_371_nl, nor_16_nl);
  assign and_1073_nl = fsm_output & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_read_1_for_mux_nl = MUX_v_8_2_2(input_read_addrs_sva_1_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4,
      and_1073_nl);
  assign or_829_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_5);
  assign nor_373_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ or_tmp_85));
  assign mux_75_nl = MUX_s_1_2_2(or_829_nl, nor_373_nl, rva_in_reg_rw_sva_st_1_5);
  assign nor_379_nl = ~((~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]!=4'b0110) | (~ reg_rva_in_PopNB_mioi_iswt0_cse));
  assign nor_380_nl = ~(nor_374_cse | reg_rva_in_reg_rw_sva_st_1_1_cse | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1));
  assign mux_77_nl = MUX_s_1_2_2(nor_379_nl, nor_380_nl, while_stage_0_3);
  assign nor_381_nl = ~((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | reg_rva_in_reg_rw_sva_2_cse | (~(accum_vector_operator_1_for_asn_73_itm_1
      | nor_375_cse)));
  assign mux_78_nl = MUX_s_1_2_2(mux_77_nl, nor_381_nl, while_stage_0_4);
  assign nor_382_nl = ~((~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1
      | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_371_itm_1 | accum_vector_operator_1_for_asn_73_itm_2))
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | rva_in_reg_rw_sva_3);
  assign mux_79_nl = MUX_s_1_2_2(mux_78_nl, nor_382_nl, while_stage_0_5);
  assign nor_383_nl = ~((~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 | rva_in_reg_rw_sva_st_1_4))
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | rva_in_reg_rw_sva_4);
  assign mux_80_nl = MUX_s_1_2_2(mux_79_nl, nor_383_nl, while_stage_0_6);
  assign mux_81_nl = MUX_s_1_2_2(mux_80_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5,
      while_stage_0_7);
  assign and_667_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign nor_499_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_234_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[15:8]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_234_nl);
  assign mux_82_nl = MUX_s_1_2_2((~ or_tmp_36), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_91_nl = MUX_s_1_2_2(and_dcpl_323, or_tmp_8, weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]);
  assign while_if_while_if_and_2_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:0])
      & ({{14{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & ({{14{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
  assign or_512_nl = or_dcpl_146 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) |
      (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | or_dcpl_305;
  assign and_748_nl = (and_747_cse | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp)
      & PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign or_334_nl = and_749_cse | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp;
  assign mux_93_nl = MUX_s_1_2_2(and_748_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      or_334_nl);
  assign mux_94_nl = MUX_s_1_2_2(mux_93_nl, (~ or_tmp_108), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1
      & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2,
      pe_manager_base_weight_sva_mx3_0, PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2,
      (pe_manager_base_weight_sva_mx2[8]), PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign mux_96_nl = MUX_s_1_2_2(not_tmp_248, or_tmp_112, weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]);
  assign mux_97_nl = MUX_s_1_2_2(not_tmp_248, or_tmp_112, weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl =
      (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[2])
      & PECore_DecodeAxiRead_switch_lp_nor_2_cse;
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl = MUX_s_1_2_2(pe_config_is_valid_sva,
      pe_manager_zero_active_sva, and_315_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl = MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1,
      (pe_manager_num_input_sva[0]), and_315_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl = MUX_v_4_2_2(pe_config_num_manager_sva,
      (pe_manager_base_bias_sva[3:0]), and_315_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl = MUX_v_7_2_2((pe_config_num_output_sva[6:0]),
      (pe_manager_base_bias_sva[14:8]), and_315_cse);
  assign mux1h_3_nl = MUX1HOT_v_4_7_2((rva_out_reg_data_55_48_sva_dfm_1_5[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_7_4,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1[7:4]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[15:12]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[15:12]),
      weight_port_read_out_data_0_1_sva_mx0_7_4, {and_1006_cse , and_1007_cse , and_1008_cse
      , and_1009_cse , and_1010_cse , and_1011_cse , nor_506_cse});
  assign not_2368_nl = ~ or_dcpl;
  assign mux1h_15_nl = MUX1HOT_v_4_7_2((rva_out_reg_data_55_48_sva_dfm_1_5[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_3_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1[3:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[11:8]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[11:8]),
      weight_port_read_out_data_0_1_sva_mx0_3_0, {and_1006_cse , and_1007_cse , and_1008_cse
      , and_1009_cse , and_1010_cse , and_1011_cse , nor_506_cse});
  assign not_2277_nl = ~ or_dcpl;
  assign mux1h_13_nl = MUX1HOT_v_7_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[30:24]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[30:24]),
      weight_port_read_out_data_0_3_sva_mx0_6_0, {and_1006_cse , and_1007_cse , and_1008_cse
      , and_1009_cse , and_1010_cse , and_1011_cse , nor_506_cse});
  assign not_2366_nl = ~ or_dcpl;
  assign mux1h_4_nl = MUX1HOT_s_1_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[31]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[31]),
      weight_port_read_out_data_0_3_sva_mx0_7, {and_1006_cse , and_1007_cse , and_1008_cse
      , and_1009_cse , and_1010_cse , and_1011_cse , nor_506_cse});
  assign mux1h_5_nl = MUX1HOT_s_1_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[23]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[23]),
      weight_port_read_out_data_0_2_sva_mx0_7, {and_1022_ssc , and_1023_cse , and_1024_cse
      , and_1025_cse , and_1026_cse , and_1027_cse , nor_508_cse});
  assign mux1h_14_nl = MUX1HOT_v_7_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[22:16]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[22:16]),
      weight_port_read_out_data_0_2_sva_mx0_6_0, {and_1022_ssc , and_1023_cse , and_1024_cse
      , and_1025_cse , and_1026_cse , and_1027_cse , nor_508_cse});
  assign not_2367_nl = ~ or_dcpl_329;
  assign weight_mem_banks_load_store_for_else_mux1h_3_nl = MUX1HOT_v_4_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[15:12]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[15:12]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[15:12]),
      {and_dcpl_631 , and_dcpl_633 , and_dcpl_634});
  assign not_2269_nl = ~ or_dcpl_331;
  assign weight_mem_banks_load_store_for_else_mux1h_87_nl = MUX1HOT_v_4_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[11:8]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[11:8]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[11:8]),
      rva_out_reg_data_39_36_sva_dfm_1_4, {and_dcpl_631 , and_dcpl_633 , and_dcpl_634
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2270_nl = ~ or_dcpl_331;
  assign weight_mem_banks_load_store_for_else_mux1h_76_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[31]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[31]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[31]),
      {and_dcpl_631 , and_dcpl_633 , and_dcpl_634});
  assign weight_mem_banks_load_store_for_else_mux1h_88_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[30:24]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[30:24]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[30:24]),
      rva_out_reg_data_62_56_sva_dfm_1_4, {and_dcpl_631 , and_dcpl_633 , and_dcpl_634
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2272_nl = ~ or_dcpl_331;
  assign weight_mem_banks_load_store_for_else_mux1h_81_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[23]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[23]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[23]),
      {and_dcpl_631 , and_dcpl_633 , and_dcpl_634});
  assign weight_mem_banks_load_store_for_else_mux1h_89_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[22:16]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[22:16]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[22:16]),
      rva_out_reg_data_46_40_sva_dfm_1_4, {and_dcpl_631 , and_dcpl_633 , and_dcpl_634
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2274_nl = ~ or_dcpl_331;
  assign weight_mem_banks_load_store_for_else_mux1h_86_nl = MUX1HOT_v_4_5_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[7:4]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[7:4]), (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[7:4]),
      (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[7:4]), (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[7:4]),
      {and_652_ssc , and_653_ssc , and_655_ssc , and_658_ssc , and_661_ssc});
  assign weight_mem_banks_load_store_for_else_or_nl = MUX_v_4_2_2(weight_mem_banks_load_store_for_else_mux1h_86_nl,
      4'b1111, and_651_ssc);
  assign mux_415_nl = MUX_v_4_2_2(weight_mem_banks_load_store_for_else_or_nl, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[7:4]),
      or_dcpl_334);
  assign not_2275_nl = ~ and_dcpl_721;
  assign and_662_nl = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign weight_mem_banks_load_store_for_else_mux1h_90_nl = MUX1HOT_v_4_6_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[3:0]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[3:0]), (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[3:0]),
      (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[3:0]), (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[3:0]),
      rva_out_reg_data_35_32_sva_dfm_1_4, {and_652_ssc , and_653_ssc , and_655_ssc
      , and_658_ssc , and_661_ssc , and_662_nl});
  assign weight_mem_banks_load_store_for_else_or_1_nl = MUX_v_4_2_2(weight_mem_banks_load_store_for_else_mux1h_90_nl,
      4'b1111, and_651_ssc);
  assign mux_416_nl = MUX_v_4_2_2(weight_mem_banks_load_store_for_else_or_1_nl, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[3:0]),
      or_dcpl_334);
  assign not_2276_nl = ~ and_dcpl_721;
  assign and_1544_nl = or_931_cse & mux_tmp_512;
  assign and_1543_nl = or_928_cse & mux_tmp_512;
  assign mux_545_nl = MUX_s_1_2_2(and_1544_nl, and_1543_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_1549_nl = or_931_cse & mux_tmp_514;
  assign and_1548_nl = or_928_cse & mux_tmp_514;
  assign mux_547_nl = MUX_s_1_2_2(and_1549_nl, and_1548_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[87:84]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_240_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_134_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[83:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_240_nl);

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_9_2;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [8:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_8_2;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [7:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    result = result | (input_5 & {11{sel[5]}});
    result = result | (input_6 & {11{sel[6]}});
    result = result | (input_7 & {11{sel[7]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function automatic [127:0] MUX1HOT_v_128_3_2;
    input [127:0] input_2;
    input [127:0] input_1;
    input [127:0] input_0;
    input [2:0] sel;
    reg [127:0] result;
  begin
    result = input_0 & {128{sel[0]}};
    result = result | (input_1 & {128{sel[1]}});
    result = result | (input_2 & {128{sel[2]}});
    MUX1HOT_v_128_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_6_2;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [5:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    MUX1HOT_v_4_6_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_7_2;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [6:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    MUX1HOT_v_4_7_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_9_2;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [8:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    MUX1HOT_v_4_9_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_7_2;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [6:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    result = result | (input_6 & {7{sel[6]}});
    MUX1HOT_v_7_7_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_9_2;
    input [6:0] input_8;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [8:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    result = result | (input_6 & {7{sel[6]}});
    result = result | (input_7 & {7{sel[7]}});
    result = result | (input_8 & {7{sel[8]}});
    MUX1HOT_v_7_9_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_7_2;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [6:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    MUX1HOT_v_8_7_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_8_2;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [7:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    MUX1HOT_v_8_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_9_2;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [8:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    result = result | (input_8 & {8{sel[8]}});
    MUX1HOT_v_8_9_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_8_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input [2:0] sel;
    reg  result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_s_1_8_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_8_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [10:0] input_2;
    input [10:0] input_3;
    input [10:0] input_4;
    input [10:0] input_5;
    input [10:0] input_6;
    input [10:0] input_7;
    input [2:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_11_8_2 = result;
  end
  endfunction


  function automatic [119:0] MUX_v_120_2_2;
    input [119:0] input_0;
    input [119:0] input_1;
    input  sel;
    reg [119:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_120_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_256_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [127:0] input_2;
    input [127:0] input_3;
    input [127:0] input_4;
    input [127:0] input_5;
    input [127:0] input_6;
    input [127:0] input_7;
    input [127:0] input_8;
    input [127:0] input_9;
    input [127:0] input_10;
    input [127:0] input_11;
    input [127:0] input_12;
    input [127:0] input_13;
    input [127:0] input_14;
    input [127:0] input_15;
    input [127:0] input_16;
    input [127:0] input_17;
    input [127:0] input_18;
    input [127:0] input_19;
    input [127:0] input_20;
    input [127:0] input_21;
    input [127:0] input_22;
    input [127:0] input_23;
    input [127:0] input_24;
    input [127:0] input_25;
    input [127:0] input_26;
    input [127:0] input_27;
    input [127:0] input_28;
    input [127:0] input_29;
    input [127:0] input_30;
    input [127:0] input_31;
    input [127:0] input_32;
    input [127:0] input_33;
    input [127:0] input_34;
    input [127:0] input_35;
    input [127:0] input_36;
    input [127:0] input_37;
    input [127:0] input_38;
    input [127:0] input_39;
    input [127:0] input_40;
    input [127:0] input_41;
    input [127:0] input_42;
    input [127:0] input_43;
    input [127:0] input_44;
    input [127:0] input_45;
    input [127:0] input_46;
    input [127:0] input_47;
    input [127:0] input_48;
    input [127:0] input_49;
    input [127:0] input_50;
    input [127:0] input_51;
    input [127:0] input_52;
    input [127:0] input_53;
    input [127:0] input_54;
    input [127:0] input_55;
    input [127:0] input_56;
    input [127:0] input_57;
    input [127:0] input_58;
    input [127:0] input_59;
    input [127:0] input_60;
    input [127:0] input_61;
    input [127:0] input_62;
    input [127:0] input_63;
    input [127:0] input_64;
    input [127:0] input_65;
    input [127:0] input_66;
    input [127:0] input_67;
    input [127:0] input_68;
    input [127:0] input_69;
    input [127:0] input_70;
    input [127:0] input_71;
    input [127:0] input_72;
    input [127:0] input_73;
    input [127:0] input_74;
    input [127:0] input_75;
    input [127:0] input_76;
    input [127:0] input_77;
    input [127:0] input_78;
    input [127:0] input_79;
    input [127:0] input_80;
    input [127:0] input_81;
    input [127:0] input_82;
    input [127:0] input_83;
    input [127:0] input_84;
    input [127:0] input_85;
    input [127:0] input_86;
    input [127:0] input_87;
    input [127:0] input_88;
    input [127:0] input_89;
    input [127:0] input_90;
    input [127:0] input_91;
    input [127:0] input_92;
    input [127:0] input_93;
    input [127:0] input_94;
    input [127:0] input_95;
    input [127:0] input_96;
    input [127:0] input_97;
    input [127:0] input_98;
    input [127:0] input_99;
    input [127:0] input_100;
    input [127:0] input_101;
    input [127:0] input_102;
    input [127:0] input_103;
    input [127:0] input_104;
    input [127:0] input_105;
    input [127:0] input_106;
    input [127:0] input_107;
    input [127:0] input_108;
    input [127:0] input_109;
    input [127:0] input_110;
    input [127:0] input_111;
    input [127:0] input_112;
    input [127:0] input_113;
    input [127:0] input_114;
    input [127:0] input_115;
    input [127:0] input_116;
    input [127:0] input_117;
    input [127:0] input_118;
    input [127:0] input_119;
    input [127:0] input_120;
    input [127:0] input_121;
    input [127:0] input_122;
    input [127:0] input_123;
    input [127:0] input_124;
    input [127:0] input_125;
    input [127:0] input_126;
    input [127:0] input_127;
    input [127:0] input_128;
    input [127:0] input_129;
    input [127:0] input_130;
    input [127:0] input_131;
    input [127:0] input_132;
    input [127:0] input_133;
    input [127:0] input_134;
    input [127:0] input_135;
    input [127:0] input_136;
    input [127:0] input_137;
    input [127:0] input_138;
    input [127:0] input_139;
    input [127:0] input_140;
    input [127:0] input_141;
    input [127:0] input_142;
    input [127:0] input_143;
    input [127:0] input_144;
    input [127:0] input_145;
    input [127:0] input_146;
    input [127:0] input_147;
    input [127:0] input_148;
    input [127:0] input_149;
    input [127:0] input_150;
    input [127:0] input_151;
    input [127:0] input_152;
    input [127:0] input_153;
    input [127:0] input_154;
    input [127:0] input_155;
    input [127:0] input_156;
    input [127:0] input_157;
    input [127:0] input_158;
    input [127:0] input_159;
    input [127:0] input_160;
    input [127:0] input_161;
    input [127:0] input_162;
    input [127:0] input_163;
    input [127:0] input_164;
    input [127:0] input_165;
    input [127:0] input_166;
    input [127:0] input_167;
    input [127:0] input_168;
    input [127:0] input_169;
    input [127:0] input_170;
    input [127:0] input_171;
    input [127:0] input_172;
    input [127:0] input_173;
    input [127:0] input_174;
    input [127:0] input_175;
    input [127:0] input_176;
    input [127:0] input_177;
    input [127:0] input_178;
    input [127:0] input_179;
    input [127:0] input_180;
    input [127:0] input_181;
    input [127:0] input_182;
    input [127:0] input_183;
    input [127:0] input_184;
    input [127:0] input_185;
    input [127:0] input_186;
    input [127:0] input_187;
    input [127:0] input_188;
    input [127:0] input_189;
    input [127:0] input_190;
    input [127:0] input_191;
    input [127:0] input_192;
    input [127:0] input_193;
    input [127:0] input_194;
    input [127:0] input_195;
    input [127:0] input_196;
    input [127:0] input_197;
    input [127:0] input_198;
    input [127:0] input_199;
    input [127:0] input_200;
    input [127:0] input_201;
    input [127:0] input_202;
    input [127:0] input_203;
    input [127:0] input_204;
    input [127:0] input_205;
    input [127:0] input_206;
    input [127:0] input_207;
    input [127:0] input_208;
    input [127:0] input_209;
    input [127:0] input_210;
    input [127:0] input_211;
    input [127:0] input_212;
    input [127:0] input_213;
    input [127:0] input_214;
    input [127:0] input_215;
    input [127:0] input_216;
    input [127:0] input_217;
    input [127:0] input_218;
    input [127:0] input_219;
    input [127:0] input_220;
    input [127:0] input_221;
    input [127:0] input_222;
    input [127:0] input_223;
    input [127:0] input_224;
    input [127:0] input_225;
    input [127:0] input_226;
    input [127:0] input_227;
    input [127:0] input_228;
    input [127:0] input_229;
    input [127:0] input_230;
    input [127:0] input_231;
    input [127:0] input_232;
    input [127:0] input_233;
    input [127:0] input_234;
    input [127:0] input_235;
    input [127:0] input_236;
    input [127:0] input_237;
    input [127:0] input_238;
    input [127:0] input_239;
    input [127:0] input_240;
    input [127:0] input_241;
    input [127:0] input_242;
    input [127:0] input_243;
    input [127:0] input_244;
    input [127:0] input_245;
    input [127:0] input_246;
    input [127:0] input_247;
    input [127:0] input_248;
    input [127:0] input_249;
    input [127:0] input_250;
    input [127:0] input_251;
    input [127:0] input_252;
    input [127:0] input_253;
    input [127:0] input_254;
    input [127:0] input_255;
    input [7:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      8'b00000000 : begin
        result = input_0;
      end
      8'b00000001 : begin
        result = input_1;
      end
      8'b00000010 : begin
        result = input_2;
      end
      8'b00000011 : begin
        result = input_3;
      end
      8'b00000100 : begin
        result = input_4;
      end
      8'b00000101 : begin
        result = input_5;
      end
      8'b00000110 : begin
        result = input_6;
      end
      8'b00000111 : begin
        result = input_7;
      end
      8'b00001000 : begin
        result = input_8;
      end
      8'b00001001 : begin
        result = input_9;
      end
      8'b00001010 : begin
        result = input_10;
      end
      8'b00001011 : begin
        result = input_11;
      end
      8'b00001100 : begin
        result = input_12;
      end
      8'b00001101 : begin
        result = input_13;
      end
      8'b00001110 : begin
        result = input_14;
      end
      8'b00001111 : begin
        result = input_15;
      end
      8'b00010000 : begin
        result = input_16;
      end
      8'b00010001 : begin
        result = input_17;
      end
      8'b00010010 : begin
        result = input_18;
      end
      8'b00010011 : begin
        result = input_19;
      end
      8'b00010100 : begin
        result = input_20;
      end
      8'b00010101 : begin
        result = input_21;
      end
      8'b00010110 : begin
        result = input_22;
      end
      8'b00010111 : begin
        result = input_23;
      end
      8'b00011000 : begin
        result = input_24;
      end
      8'b00011001 : begin
        result = input_25;
      end
      8'b00011010 : begin
        result = input_26;
      end
      8'b00011011 : begin
        result = input_27;
      end
      8'b00011100 : begin
        result = input_28;
      end
      8'b00011101 : begin
        result = input_29;
      end
      8'b00011110 : begin
        result = input_30;
      end
      8'b00011111 : begin
        result = input_31;
      end
      8'b00100000 : begin
        result = input_32;
      end
      8'b00100001 : begin
        result = input_33;
      end
      8'b00100010 : begin
        result = input_34;
      end
      8'b00100011 : begin
        result = input_35;
      end
      8'b00100100 : begin
        result = input_36;
      end
      8'b00100101 : begin
        result = input_37;
      end
      8'b00100110 : begin
        result = input_38;
      end
      8'b00100111 : begin
        result = input_39;
      end
      8'b00101000 : begin
        result = input_40;
      end
      8'b00101001 : begin
        result = input_41;
      end
      8'b00101010 : begin
        result = input_42;
      end
      8'b00101011 : begin
        result = input_43;
      end
      8'b00101100 : begin
        result = input_44;
      end
      8'b00101101 : begin
        result = input_45;
      end
      8'b00101110 : begin
        result = input_46;
      end
      8'b00101111 : begin
        result = input_47;
      end
      8'b00110000 : begin
        result = input_48;
      end
      8'b00110001 : begin
        result = input_49;
      end
      8'b00110010 : begin
        result = input_50;
      end
      8'b00110011 : begin
        result = input_51;
      end
      8'b00110100 : begin
        result = input_52;
      end
      8'b00110101 : begin
        result = input_53;
      end
      8'b00110110 : begin
        result = input_54;
      end
      8'b00110111 : begin
        result = input_55;
      end
      8'b00111000 : begin
        result = input_56;
      end
      8'b00111001 : begin
        result = input_57;
      end
      8'b00111010 : begin
        result = input_58;
      end
      8'b00111011 : begin
        result = input_59;
      end
      8'b00111100 : begin
        result = input_60;
      end
      8'b00111101 : begin
        result = input_61;
      end
      8'b00111110 : begin
        result = input_62;
      end
      8'b00111111 : begin
        result = input_63;
      end
      8'b01000000 : begin
        result = input_64;
      end
      8'b01000001 : begin
        result = input_65;
      end
      8'b01000010 : begin
        result = input_66;
      end
      8'b01000011 : begin
        result = input_67;
      end
      8'b01000100 : begin
        result = input_68;
      end
      8'b01000101 : begin
        result = input_69;
      end
      8'b01000110 : begin
        result = input_70;
      end
      8'b01000111 : begin
        result = input_71;
      end
      8'b01001000 : begin
        result = input_72;
      end
      8'b01001001 : begin
        result = input_73;
      end
      8'b01001010 : begin
        result = input_74;
      end
      8'b01001011 : begin
        result = input_75;
      end
      8'b01001100 : begin
        result = input_76;
      end
      8'b01001101 : begin
        result = input_77;
      end
      8'b01001110 : begin
        result = input_78;
      end
      8'b01001111 : begin
        result = input_79;
      end
      8'b01010000 : begin
        result = input_80;
      end
      8'b01010001 : begin
        result = input_81;
      end
      8'b01010010 : begin
        result = input_82;
      end
      8'b01010011 : begin
        result = input_83;
      end
      8'b01010100 : begin
        result = input_84;
      end
      8'b01010101 : begin
        result = input_85;
      end
      8'b01010110 : begin
        result = input_86;
      end
      8'b01010111 : begin
        result = input_87;
      end
      8'b01011000 : begin
        result = input_88;
      end
      8'b01011001 : begin
        result = input_89;
      end
      8'b01011010 : begin
        result = input_90;
      end
      8'b01011011 : begin
        result = input_91;
      end
      8'b01011100 : begin
        result = input_92;
      end
      8'b01011101 : begin
        result = input_93;
      end
      8'b01011110 : begin
        result = input_94;
      end
      8'b01011111 : begin
        result = input_95;
      end
      8'b01100000 : begin
        result = input_96;
      end
      8'b01100001 : begin
        result = input_97;
      end
      8'b01100010 : begin
        result = input_98;
      end
      8'b01100011 : begin
        result = input_99;
      end
      8'b01100100 : begin
        result = input_100;
      end
      8'b01100101 : begin
        result = input_101;
      end
      8'b01100110 : begin
        result = input_102;
      end
      8'b01100111 : begin
        result = input_103;
      end
      8'b01101000 : begin
        result = input_104;
      end
      8'b01101001 : begin
        result = input_105;
      end
      8'b01101010 : begin
        result = input_106;
      end
      8'b01101011 : begin
        result = input_107;
      end
      8'b01101100 : begin
        result = input_108;
      end
      8'b01101101 : begin
        result = input_109;
      end
      8'b01101110 : begin
        result = input_110;
      end
      8'b01101111 : begin
        result = input_111;
      end
      8'b01110000 : begin
        result = input_112;
      end
      8'b01110001 : begin
        result = input_113;
      end
      8'b01110010 : begin
        result = input_114;
      end
      8'b01110011 : begin
        result = input_115;
      end
      8'b01110100 : begin
        result = input_116;
      end
      8'b01110101 : begin
        result = input_117;
      end
      8'b01110110 : begin
        result = input_118;
      end
      8'b01110111 : begin
        result = input_119;
      end
      8'b01111000 : begin
        result = input_120;
      end
      8'b01111001 : begin
        result = input_121;
      end
      8'b01111010 : begin
        result = input_122;
      end
      8'b01111011 : begin
        result = input_123;
      end
      8'b01111100 : begin
        result = input_124;
      end
      8'b01111101 : begin
        result = input_125;
      end
      8'b01111110 : begin
        result = input_126;
      end
      8'b01111111 : begin
        result = input_127;
      end
      8'b10000000 : begin
        result = input_128;
      end
      8'b10000001 : begin
        result = input_129;
      end
      8'b10000010 : begin
        result = input_130;
      end
      8'b10000011 : begin
        result = input_131;
      end
      8'b10000100 : begin
        result = input_132;
      end
      8'b10000101 : begin
        result = input_133;
      end
      8'b10000110 : begin
        result = input_134;
      end
      8'b10000111 : begin
        result = input_135;
      end
      8'b10001000 : begin
        result = input_136;
      end
      8'b10001001 : begin
        result = input_137;
      end
      8'b10001010 : begin
        result = input_138;
      end
      8'b10001011 : begin
        result = input_139;
      end
      8'b10001100 : begin
        result = input_140;
      end
      8'b10001101 : begin
        result = input_141;
      end
      8'b10001110 : begin
        result = input_142;
      end
      8'b10001111 : begin
        result = input_143;
      end
      8'b10010000 : begin
        result = input_144;
      end
      8'b10010001 : begin
        result = input_145;
      end
      8'b10010010 : begin
        result = input_146;
      end
      8'b10010011 : begin
        result = input_147;
      end
      8'b10010100 : begin
        result = input_148;
      end
      8'b10010101 : begin
        result = input_149;
      end
      8'b10010110 : begin
        result = input_150;
      end
      8'b10010111 : begin
        result = input_151;
      end
      8'b10011000 : begin
        result = input_152;
      end
      8'b10011001 : begin
        result = input_153;
      end
      8'b10011010 : begin
        result = input_154;
      end
      8'b10011011 : begin
        result = input_155;
      end
      8'b10011100 : begin
        result = input_156;
      end
      8'b10011101 : begin
        result = input_157;
      end
      8'b10011110 : begin
        result = input_158;
      end
      8'b10011111 : begin
        result = input_159;
      end
      8'b10100000 : begin
        result = input_160;
      end
      8'b10100001 : begin
        result = input_161;
      end
      8'b10100010 : begin
        result = input_162;
      end
      8'b10100011 : begin
        result = input_163;
      end
      8'b10100100 : begin
        result = input_164;
      end
      8'b10100101 : begin
        result = input_165;
      end
      8'b10100110 : begin
        result = input_166;
      end
      8'b10100111 : begin
        result = input_167;
      end
      8'b10101000 : begin
        result = input_168;
      end
      8'b10101001 : begin
        result = input_169;
      end
      8'b10101010 : begin
        result = input_170;
      end
      8'b10101011 : begin
        result = input_171;
      end
      8'b10101100 : begin
        result = input_172;
      end
      8'b10101101 : begin
        result = input_173;
      end
      8'b10101110 : begin
        result = input_174;
      end
      8'b10101111 : begin
        result = input_175;
      end
      8'b10110000 : begin
        result = input_176;
      end
      8'b10110001 : begin
        result = input_177;
      end
      8'b10110010 : begin
        result = input_178;
      end
      8'b10110011 : begin
        result = input_179;
      end
      8'b10110100 : begin
        result = input_180;
      end
      8'b10110101 : begin
        result = input_181;
      end
      8'b10110110 : begin
        result = input_182;
      end
      8'b10110111 : begin
        result = input_183;
      end
      8'b10111000 : begin
        result = input_184;
      end
      8'b10111001 : begin
        result = input_185;
      end
      8'b10111010 : begin
        result = input_186;
      end
      8'b10111011 : begin
        result = input_187;
      end
      8'b10111100 : begin
        result = input_188;
      end
      8'b10111101 : begin
        result = input_189;
      end
      8'b10111110 : begin
        result = input_190;
      end
      8'b10111111 : begin
        result = input_191;
      end
      8'b11000000 : begin
        result = input_192;
      end
      8'b11000001 : begin
        result = input_193;
      end
      8'b11000010 : begin
        result = input_194;
      end
      8'b11000011 : begin
        result = input_195;
      end
      8'b11000100 : begin
        result = input_196;
      end
      8'b11000101 : begin
        result = input_197;
      end
      8'b11000110 : begin
        result = input_198;
      end
      8'b11000111 : begin
        result = input_199;
      end
      8'b11001000 : begin
        result = input_200;
      end
      8'b11001001 : begin
        result = input_201;
      end
      8'b11001010 : begin
        result = input_202;
      end
      8'b11001011 : begin
        result = input_203;
      end
      8'b11001100 : begin
        result = input_204;
      end
      8'b11001101 : begin
        result = input_205;
      end
      8'b11001110 : begin
        result = input_206;
      end
      8'b11001111 : begin
        result = input_207;
      end
      8'b11010000 : begin
        result = input_208;
      end
      8'b11010001 : begin
        result = input_209;
      end
      8'b11010010 : begin
        result = input_210;
      end
      8'b11010011 : begin
        result = input_211;
      end
      8'b11010100 : begin
        result = input_212;
      end
      8'b11010101 : begin
        result = input_213;
      end
      8'b11010110 : begin
        result = input_214;
      end
      8'b11010111 : begin
        result = input_215;
      end
      8'b11011000 : begin
        result = input_216;
      end
      8'b11011001 : begin
        result = input_217;
      end
      8'b11011010 : begin
        result = input_218;
      end
      8'b11011011 : begin
        result = input_219;
      end
      8'b11011100 : begin
        result = input_220;
      end
      8'b11011101 : begin
        result = input_221;
      end
      8'b11011110 : begin
        result = input_222;
      end
      8'b11011111 : begin
        result = input_223;
      end
      8'b11100000 : begin
        result = input_224;
      end
      8'b11100001 : begin
        result = input_225;
      end
      8'b11100010 : begin
        result = input_226;
      end
      8'b11100011 : begin
        result = input_227;
      end
      8'b11100100 : begin
        result = input_228;
      end
      8'b11100101 : begin
        result = input_229;
      end
      8'b11100110 : begin
        result = input_230;
      end
      8'b11100111 : begin
        result = input_231;
      end
      8'b11101000 : begin
        result = input_232;
      end
      8'b11101001 : begin
        result = input_233;
      end
      8'b11101010 : begin
        result = input_234;
      end
      8'b11101011 : begin
        result = input_235;
      end
      8'b11101100 : begin
        result = input_236;
      end
      8'b11101101 : begin
        result = input_237;
      end
      8'b11101110 : begin
        result = input_238;
      end
      8'b11101111 : begin
        result = input_239;
      end
      8'b11110000 : begin
        result = input_240;
      end
      8'b11110001 : begin
        result = input_241;
      end
      8'b11110010 : begin
        result = input_242;
      end
      8'b11110011 : begin
        result = input_243;
      end
      8'b11110100 : begin
        result = input_244;
      end
      8'b11110101 : begin
        result = input_245;
      end
      8'b11110110 : begin
        result = input_246;
      end
      8'b11110111 : begin
        result = input_247;
      end
      8'b11111000 : begin
        result = input_248;
      end
      8'b11111001 : begin
        result = input_249;
      end
      8'b11111010 : begin
        result = input_250;
      end
      8'b11111011 : begin
        result = input_251;
      end
      8'b11111100 : begin
        result = input_252;
      end
      8'b11111101 : begin
        result = input_253;
      end
      8'b11111110 : begin
        result = input_254;
      end
      default : begin
        result = input_255;
      end
    endcase
    MUX_v_128_256_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input  sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input  sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [27:0] MUX_v_28_2_2;
    input [27:0] input_0;
    input [27:0] input_1;
    input  sel;
    reg [27:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_28_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_8_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [1:0] input_2;
    input [1:0] input_3;
    input [1:0] input_4;
    input [1:0] input_5;
    input [1:0] input_6;
    input [1:0] input_7;
    input [2:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_2_8_2 = result;
  end
  endfunction


  function automatic [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input  sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_8_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [2:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_4_8_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_8_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [5:0] input_2;
    input [5:0] input_3;
    input [5:0] input_4;
    input [5:0] input_5;
    input [5:0] input_6;
    input [5:0] input_7;
    input [2:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_6_8_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_8_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [6:0] input_2;
    input [6:0] input_3;
    input [6:0] input_4;
    input [6:0] input_5;
    input [6:0] input_6;
    input [6:0] input_7;
    input [2:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_7_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [10:0] signext_11_1;
    input  vector;
  begin
    signext_11_1= {{10{vector}}, vector};
  end
  endfunction


  function automatic [255:0] signext_256_252;
    input [251:0] vector;
  begin
    signext_256_252= {{4{vector[251]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [31:0] signext_32_28;
    input [27:0] vector;
  begin
    signext_32_28= {{4{vector[27]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input  vector;
  begin
    signext_3_1= {{2{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input  vector;
  begin
    signext_4_1= {{3{vector}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input  vector;
  begin
    signext_7_1= {{6{vector}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore
// ------------------------------------------------------------------


module PECore (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [137:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  wire [7:0] ProductSum_for_acc_20_cmp_a;
  wire ProductSum_for_acc_20_cmp_load;
  wire ProductSum_for_acc_20_cmp_en;
  wire [30:0] ProductSum_for_acc_20_cmp_z;
  wire [7:0] ProductSum_for_acc_19_cmp_a0;
  wire [7:0] ProductSum_for_acc_19_cmp_b0;
  wire [7:0] ProductSum_for_acc_19_cmp_c0;
  wire ProductSum_for_acc_19_cmp_en;
  wire [30:0] ProductSum_for_acc_19_cmp_z;
  wire [7:0] ProductSum_for_acc_18_cmp_a0;
  wire [7:0] ProductSum_for_acc_18_cmp_b0;
  wire [7:0] ProductSum_for_acc_18_cmp_c0;
  wire [30:0] ProductSum_for_acc_18_cmp_z;
  wire [7:0] ProductSum_for_acc_17_cmp_a0;
  wire [7:0] ProductSum_for_acc_17_cmp_b0;
  wire [7:0] ProductSum_for_acc_17_cmp_c0;
  wire [30:0] ProductSum_for_acc_17_cmp_z;
  wire [7:0] ProductSum_for_acc_16_cmp_a0;
  wire [7:0] ProductSum_for_acc_16_cmp_b0;
  wire [7:0] ProductSum_for_acc_16_cmp_c0;
  wire [30:0] ProductSum_for_acc_16_cmp_z;
  wire [7:0] ProductSum_for_acc_15_cmp_a0;
  wire [7:0] ProductSum_for_acc_15_cmp_b0;
  wire [7:0] ProductSum_for_acc_15_cmp_c0;
  wire [30:0] ProductSum_for_acc_15_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_a;
  wire PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_load;
  wire [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_a;
  wire PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_load;
  wire [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_a;
  wire [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_a;
  wire PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_load;
  wire [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_a;
  wire [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_a;
  wire PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_load;
  wire [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_a;
  wire PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_load;
  wire [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [30:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr;
  wire [7:0] ProductSum_for_acc_20_cmp_b_iff;
  wire ProductSum_for_acc_20_cmp_datavalid_iff;
  wire [7:0] ProductSum_for_acc_19_cmp_a1_iff;
  wire [7:0] ProductSum_for_acc_19_cmp_b1_iff;
  wire [7:0] ProductSum_for_acc_19_cmp_c1_iff;
  wire ProductSum_for_acc_19_cmp_load_iff;
  wire ProductSum_for_acc_19_cmp_datavalid_iff;
  wire [7:0] ProductSum_for_acc_18_cmp_a1_iff;
  wire [7:0] ProductSum_for_acc_18_cmp_b1_iff;
  wire [7:0] ProductSum_for_acc_18_cmp_c1_iff;
  wire [7:0] ProductSum_for_acc_17_cmp_a1_iff;
  wire [7:0] ProductSum_for_acc_17_cmp_b1_iff;
  wire [7:0] ProductSum_for_acc_17_cmp_c1_iff;
  wire [7:0] ProductSum_for_acc_16_cmp_a1_iff;
  wire [7:0] ProductSum_for_acc_16_cmp_b1_iff;
  wire [7:0] ProductSum_for_acc_16_cmp_c1_iff;
  wire [7:0] ProductSum_for_acc_15_cmp_a1_iff;
  wire [7:0] ProductSum_for_acc_15_cmp_b1_iff;
  wire [7:0] ProductSum_for_acc_15_cmp_c1_iff;
  wire PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_iff;
  wire PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_iff;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_b_iff;
  wire PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_iff;
  wire PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_iff;
  wire PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_iff;
  wire PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_iff;
  wire PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd31),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd31),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_20_cmp (
      .a(ProductSum_for_acc_20_cmp_a),
      .b(ProductSum_for_acc_20_cmp_b_iff),
      .c(31'b0000000000000000000000000000000),
      .load(ProductSum_for_acc_20_cmp_load),
      .datavalid(ProductSum_for_acc_20_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_20_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_20_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_19_cmp (
      .a0(ProductSum_for_acc_19_cmp_a0),
      .a1(ProductSum_for_acc_19_cmp_a1_iff),
      .b0(ProductSum_for_acc_19_cmp_b0),
      .b1(ProductSum_for_acc_19_cmp_b1_iff),
      .c0(ProductSum_for_acc_19_cmp_c0),
      .c1(ProductSum_for_acc_19_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(ProductSum_for_acc_19_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_19_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_18_cmp (
      .a0(ProductSum_for_acc_18_cmp_a0),
      .a1(ProductSum_for_acc_18_cmp_a1_iff),
      .b0(ProductSum_for_acc_18_cmp_b0),
      .b1(ProductSum_for_acc_18_cmp_b1_iff),
      .c0(ProductSum_for_acc_18_cmp_c0),
      .c1(ProductSum_for_acc_18_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(ProductSum_for_acc_19_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_18_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_17_cmp (
      .a0(ProductSum_for_acc_17_cmp_a0),
      .a1(ProductSum_for_acc_17_cmp_a1_iff),
      .b0(ProductSum_for_acc_17_cmp_b0),
      .b1(ProductSum_for_acc_17_cmp_b1_iff),
      .c0(ProductSum_for_acc_17_cmp_c0),
      .c1(ProductSum_for_acc_17_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(ProductSum_for_acc_19_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_17_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_16_cmp (
      .a0(ProductSum_for_acc_16_cmp_a0),
      .a1(ProductSum_for_acc_16_cmp_a1_iff),
      .b0(ProductSum_for_acc_16_cmp_b0),
      .b1(ProductSum_for_acc_16_cmp_b1_iff),
      .c0(ProductSum_for_acc_16_cmp_c0),
      .c1(ProductSum_for_acc_16_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(ProductSum_for_acc_19_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_16_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_15_cmp (
      .a0(ProductSum_for_acc_15_cmp_a0),
      .a1(ProductSum_for_acc_15_cmp_a1_iff),
      .b0(ProductSum_for_acc_15_cmp_b0),
      .b1(ProductSum_for_acc_15_cmp_b1_iff),
      .c0(ProductSum_for_acc_15_cmp_c0),
      .c1(ProductSum_for_acc_15_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(ProductSum_for_acc_19_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_15_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd31),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd31),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp (
      .a(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .b(ProductSum_for_acc_20_cmp_b_iff),
      .c(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .datavalid(ProductSum_for_acc_20_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_20_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp (
      .a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .a1(ProductSum_for_acc_19_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .b1(ProductSum_for_acc_19_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .c1(ProductSum_for_acc_19_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp (
      .a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .a1(ProductSum_for_acc_18_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .b1(ProductSum_for_acc_18_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .c1(ProductSum_for_acc_18_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp (
      .a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .a1(ProductSum_for_acc_17_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .b1(ProductSum_for_acc_17_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .c1(ProductSum_for_acc_17_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_16_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_16_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_16_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_15_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_15_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_15_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd31),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd31),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp (
      .a(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .b(ProductSum_for_acc_20_cmp_b_iff),
      .c(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .datavalid(ProductSum_for_acc_20_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_20_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp (
      .a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .a1(ProductSum_for_acc_19_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .b1(ProductSum_for_acc_19_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .c1(ProductSum_for_acc_19_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp (
      .a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .a1(ProductSum_for_acc_18_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .b1(ProductSum_for_acc_18_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .c1(ProductSum_for_acc_18_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp (
      .a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .a1(ProductSum_for_acc_17_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .b1(ProductSum_for_acc_17_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .c1(ProductSum_for_acc_17_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_16_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_16_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_16_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_15_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_15_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_15_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd31),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd31),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp (
      .a(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .b(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_b_iff),
      .c(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp (
      .a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .a1(ProductSum_for_acc_19_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .b1(ProductSum_for_acc_19_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .c1(ProductSum_for_acc_19_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp (
      .a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .a1(ProductSum_for_acc_18_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .b1(ProductSum_for_acc_18_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .c1(ProductSum_for_acc_18_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp (
      .a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .a1(ProductSum_for_acc_17_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .b1(ProductSum_for_acc_17_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .c1(ProductSum_for_acc_17_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_16_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_16_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_16_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_15_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_15_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_15_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd31),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd31),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp (
      .a(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .b(ProductSum_for_acc_20_cmp_b_iff),
      .c(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .datavalid(ProductSum_for_acc_20_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_20_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp (
      .a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .a1(ProductSum_for_acc_19_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .b1(ProductSum_for_acc_19_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .c1(ProductSum_for_acc_19_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp (
      .a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .a1(ProductSum_for_acc_18_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .b1(ProductSum_for_acc_18_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .c1(ProductSum_for_acc_18_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp (
      .a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .a1(ProductSum_for_acc_17_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .b1(ProductSum_for_acc_17_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .c1(ProductSum_for_acc_17_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_16_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_16_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_16_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_15_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_15_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_15_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd31),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd31),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp (
      .a(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .b(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_b_iff),
      .c(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp (
      .a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .a1(ProductSum_for_acc_19_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .b1(ProductSum_for_acc_19_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .c1(ProductSum_for_acc_19_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp (
      .a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .a1(ProductSum_for_acc_18_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .b1(ProductSum_for_acc_18_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .c1(ProductSum_for_acc_18_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp (
      .a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .a1(ProductSum_for_acc_17_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .b1(ProductSum_for_acc_17_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .c1(ProductSum_for_acc_17_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_16_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_16_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_16_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_15_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_15_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_15_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd31),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd31),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp (
      .a(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .b(ProductSum_for_acc_20_cmp_b_iff),
      .c(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .datavalid(ProductSum_for_acc_20_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_20_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp (
      .a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .a1(ProductSum_for_acc_19_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .b1(ProductSum_for_acc_19_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .c1(ProductSum_for_acc_19_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp (
      .a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .a1(ProductSum_for_acc_18_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .b1(ProductSum_for_acc_18_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .c1(ProductSum_for_acc_18_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp (
      .a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .a1(ProductSum_for_acc_17_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .b1(ProductSum_for_acc_17_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .c1(ProductSum_for_acc_17_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_16_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_16_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_16_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_15_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_15_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_15_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd31),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd31),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp (
      .a(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .b(ProductSum_for_acc_20_cmp_b_iff),
      .c(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .datavalid(ProductSum_for_acc_20_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_20_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp (
      .a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .a1(ProductSum_for_acc_19_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .b1(ProductSum_for_acc_19_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .c1(ProductSum_for_acc_19_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp (
      .a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .a1(ProductSum_for_acc_18_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .b1(ProductSum_for_acc_18_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .c1(ProductSum_for_acc_18_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp (
      .a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .a1(ProductSum_for_acc_17_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .b1(ProductSum_for_acc_17_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .c1(ProductSum_for_acc_17_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_16_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_16_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_16_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd31),
  .signd_e(32'sd1),
  .width_z(32'sd31),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_15_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_15_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_15_cmp_c1_iff),
      .e(31'b0000000000000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .datavalid(ProductSum_for_acc_19_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_19_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_139_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_PECoreRun PECore_PECoreRun_inst (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .ProductSum_for_acc_20_cmp_a(ProductSum_for_acc_20_cmp_a),
      .ProductSum_for_acc_20_cmp_load(ProductSum_for_acc_20_cmp_load),
      .ProductSum_for_acc_20_cmp_en(ProductSum_for_acc_20_cmp_en),
      .ProductSum_for_acc_20_cmp_z(ProductSum_for_acc_20_cmp_z),
      .ProductSum_for_acc_19_cmp_a0(ProductSum_for_acc_19_cmp_a0),
      .ProductSum_for_acc_19_cmp_b0(ProductSum_for_acc_19_cmp_b0),
      .ProductSum_for_acc_19_cmp_c0(ProductSum_for_acc_19_cmp_c0),
      .ProductSum_for_acc_19_cmp_en(ProductSum_for_acc_19_cmp_en),
      .ProductSum_for_acc_19_cmp_z(ProductSum_for_acc_19_cmp_z),
      .ProductSum_for_acc_18_cmp_a0(ProductSum_for_acc_18_cmp_a0),
      .ProductSum_for_acc_18_cmp_b0(ProductSum_for_acc_18_cmp_b0),
      .ProductSum_for_acc_18_cmp_c0(ProductSum_for_acc_18_cmp_c0),
      .ProductSum_for_acc_18_cmp_z(ProductSum_for_acc_18_cmp_z),
      .ProductSum_for_acc_17_cmp_a0(ProductSum_for_acc_17_cmp_a0),
      .ProductSum_for_acc_17_cmp_b0(ProductSum_for_acc_17_cmp_b0),
      .ProductSum_for_acc_17_cmp_c0(ProductSum_for_acc_17_cmp_c0),
      .ProductSum_for_acc_17_cmp_z(ProductSum_for_acc_17_cmp_z),
      .ProductSum_for_acc_16_cmp_a0(ProductSum_for_acc_16_cmp_a0),
      .ProductSum_for_acc_16_cmp_b0(ProductSum_for_acc_16_cmp_b0),
      .ProductSum_for_acc_16_cmp_c0(ProductSum_for_acc_16_cmp_c0),
      .ProductSum_for_acc_16_cmp_z(ProductSum_for_acc_16_cmp_z),
      .ProductSum_for_acc_15_cmp_a0(ProductSum_for_acc_15_cmp_a0),
      .ProductSum_for_acc_15_cmp_b0(ProductSum_for_acc_15_cmp_b0),
      .ProductSum_for_acc_15_cmp_c0(ProductSum_for_acc_15_cmp_c0),
      .ProductSum_for_acc_15_cmp_z(ProductSum_for_acc_15_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_a(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_a(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_a(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_a(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_a(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_a(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_a(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_a),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_load),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_7_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_a0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_b0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_c0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_b0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_c0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_b0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_c0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .ProductSum_for_acc_20_cmp_b_pff(ProductSum_for_acc_20_cmp_b_iff),
      .ProductSum_for_acc_20_cmp_datavalid_pff(ProductSum_for_acc_20_cmp_datavalid_iff),
      .ProductSum_for_acc_19_cmp_a1_pff(ProductSum_for_acc_19_cmp_a1_iff),
      .ProductSum_for_acc_19_cmp_b1_pff(ProductSum_for_acc_19_cmp_b1_iff),
      .ProductSum_for_acc_19_cmp_c1_pff(ProductSum_for_acc_19_cmp_c1_iff),
      .ProductSum_for_acc_19_cmp_load_pff(ProductSum_for_acc_19_cmp_load_iff),
      .ProductSum_for_acc_19_cmp_datavalid_pff(ProductSum_for_acc_19_cmp_datavalid_iff),
      .ProductSum_for_acc_18_cmp_a1_pff(ProductSum_for_acc_18_cmp_a1_iff),
      .ProductSum_for_acc_18_cmp_b1_pff(ProductSum_for_acc_18_cmp_b1_iff),
      .ProductSum_for_acc_18_cmp_c1_pff(ProductSum_for_acc_18_cmp_c1_iff),
      .ProductSum_for_acc_17_cmp_a1_pff(ProductSum_for_acc_17_cmp_a1_iff),
      .ProductSum_for_acc_17_cmp_b1_pff(ProductSum_for_acc_17_cmp_b1_iff),
      .ProductSum_for_acc_17_cmp_c1_pff(ProductSum_for_acc_17_cmp_c1_iff),
      .ProductSum_for_acc_16_cmp_a1_pff(ProductSum_for_acc_16_cmp_a1_iff),
      .ProductSum_for_acc_16_cmp_b1_pff(ProductSum_for_acc_16_cmp_b1_iff),
      .ProductSum_for_acc_16_cmp_c1_pff(ProductSum_for_acc_16_cmp_c1_iff),
      .ProductSum_for_acc_15_cmp_a1_pff(ProductSum_for_acc_15_cmp_a1_iff),
      .ProductSum_for_acc_15_cmp_b1_pff(ProductSum_for_acc_15_cmp_b1_iff),
      .ProductSum_for_acc_15_cmp_c1_pff(ProductSum_for_acc_15_cmp_c1_iff),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_pff(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_pff(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_b_pff(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_b_iff),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_pff(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_pff(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_pff(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_7_cmp_load_iff),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_pff(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_pff(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_6_cmp_load_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff)
    );
endmodule



