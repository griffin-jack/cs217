
//------> ./GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:55:48 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_wstrb_rsc_z,
      data_rw_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [168:0] this_dat;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output [15:0] data_wstrb_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [127:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_dat[127:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_dat[151:128];
  wire [15:0] nl_data_wstrb_rsci_d;
  assign nl_data_wstrb_rsci_d = this_dat[167:152];
  wire  nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_dat[168];
  GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd128)) data_data_rsci (
      .d(nl_data_data_rsci_d[127:0]),
      .z(data_data_rsc_z)
    );
  GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd3),
  .width(32'sd16)) data_wstrb_rsci (
      .d(nl_data_wstrb_rsci_d[15:0]),
      .z(data_wstrb_rsc_z)
    );
  GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d),
      .z(data_rw_rsc_z)
    );
  GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd155),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module GBModule_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_wstrb_rsc_z,
      data_rw_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [168:0] this_dat;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output [15:0] data_wstrb_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_wstrb_rsc_z(data_wstrb_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:56:04 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_is_write_rsc_dat, m_memory_index_rsc_dat, m_vector_index_rsc_dat,
      m_timestep_index_rsc_dat, m_write_data_data_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [154:0] this_dat;
  input m_is_write_rsc_dat;
  input [1:0] m_memory_index_rsc_dat;
  input [7:0] m_vector_index_rsc_dat;
  input [15:0] m_timestep_index_rsc_dat;
  input [127:0] m_write_data_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire m_is_write_rsci_idat;
  wire [1:0] m_memory_index_rsci_idat;
  wire [7:0] m_vector_index_rsci_idat;
  wire [15:0] m_timestep_index_rsci_idat;
  wire [127:0] m_write_data_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [127:0] m_write_data_data_buf_lpi_1_dfm;
  reg [7:0] m_vector_index_buf_lpi_1_dfm;
  reg [15:0] m_timestep_index_buf_lpi_1_dfm;
  reg [1:0] m_memory_index_buf_lpi_1_dfm;
  reg m_is_write_buf_lpi_1_dfm;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd92),
  .width(32'sd1)) m_is_write_rsci (
      .dat(m_is_write_rsc_dat),
      .idat(m_is_write_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd93),
  .width(32'sd2)) m_memory_index_rsci (
      .dat(m_memory_index_rsc_dat),
      .idat(m_memory_index_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd94),
  .width(32'sd8)) m_vector_index_rsci (
      .dat(m_vector_index_rsc_dat),
      .idat(m_vector_index_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd95),
  .width(32'sd16)) m_timestep_index_rsci (
      .dat(m_timestep_index_rsc_dat),
      .idat(m_timestep_index_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd96),
  .width(32'sd128)) m_write_data_data_rsci (
      .dat(m_write_data_data_rsc_dat),
      .idat(m_write_data_data_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd151),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd158)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = {m_write_data_data_buf_lpi_1_dfm , m_vector_index_buf_lpi_1_dfm
      , m_timestep_index_buf_lpi_1_dfm , m_memory_index_buf_lpi_1_dfm , m_is_write_buf_lpi_1_dfm};
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_write_data_data_buf_lpi_1_dfm <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_write_data_data_buf_lpi_1_dfm <= m_write_data_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_vector_index_buf_lpi_1_dfm <= 8'b00000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_vector_index_buf_lpi_1_dfm <= m_vector_index_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_timestep_index_buf_lpi_1_dfm <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_timestep_index_buf_lpi_1_dfm <= m_timestep_index_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_memory_index_buf_lpi_1_dfm <= 2'b00;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_memory_index_buf_lpi_1_dfm <= m_memory_index_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_is_write_buf_lpi_1_dfm <= 1'b0;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_is_write_buf_lpi_1_dfm <= m_is_write_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module GBModule_Connections_OutBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_is_write_rsc_dat, m_memory_index_rsc_dat, m_vector_index_rsc_dat,
      m_timestep_index_rsc_dat, m_write_data_data_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [154:0] this_dat;
  input m_is_write_rsc_dat;
  input [1:0] m_memory_index_rsc_dat;
  input [7:0] m_vector_index_rsc_dat;
  input [15:0] m_timestep_index_rsc_dat;
  input [127:0] m_write_data_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_is_write_rsc_dat(m_is_write_rsc_dat),
      .m_memory_index_rsc_dat(m_memory_index_rsc_dat),
      .m_vector_index_rsc_dat(m_vector_index_rsc_dat),
      .m_timestep_index_rsc_dat(m_timestep_index_rsc_dat),
      .m_write_data_data_rsc_dat(m_write_data_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:56:07 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd98),
  .width(32'sd1)) data_rsci (
      .d(this_dat),
      .z(data_rsc_z)
    );
  GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd100),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd150),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module GBModule_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:55:58 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_read_vector_data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [127:0] this_dat;
  output [127:0] data_read_vector_data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd101),
  .width(32'sd128)) data_read_vector_data_data_rsci (
      .d(this_dat),
      .z(data_read_vector_data_data_rsc_z)
    );
  GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd103),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd149),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module GBModule_Connections_InBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_read_vector_data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [127:0] this_dat;
  output [127:0] data_read_vector_data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_InBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_read_vector_data_data_rsc_z(data_read_vector_data_data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:55:40 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [127:0] this_dat;
  reg [127:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [127:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd15),
  .width(32'sd128)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd153),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd160)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module GBModule_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [127:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module GBModule_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./GBModule_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:55:55 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module GBModule_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output this_dat;
  reg this_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  GBModule_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd148),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd157)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_rdy));
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      this_dat <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_bool_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module GBModule_Connections_OutBlocking_bool_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output this_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule_mgc_shift_br_beh_v5.v 
module GBModule_mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction

endmodule

//------> ./GBModule_mgc_shift_bl_beh_v5.v 
module GBModule_mgc_shift_bl_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> ./GBModule_mgc_shift_l_beh_v5.v 
module GBModule_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./GBModule_leading_sign_32_1_1_0.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-01
//  Generated date: Wed Feb  4 22:01:26 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_32_1_1_0
// ------------------------------------------------------------------


module GBModule_leading_sign_32_1_1_0 (
  mantissa, all_same, rtn
);
  input [31:0] mantissa;
  output all_same;
  output [4:0] rtn;


  // Interconnect Declarations
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_2;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_42_4_sdt_4;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_50_2_sdt_2;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_62_3_sdt_3;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_70_2_sdt_2;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_76_2_sdt_1;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_90_5_sdt_5;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_34_2_sdt_1;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_50_2_sdt_1;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_58_2_sdt_1;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_70_2_sdt_1;
  wire [30:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;

  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_117_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_115_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_124_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_125_nl;

  // Interconnect Declarations for Component Instantiations
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0 =
      (mantissa[30:0]) ^ (signext_31_1(~ (mantissa[31])));
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[28:27]==2'b11);
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[30:29]==2'b11);
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[26:25]==2'b11);
  assign c_h_1_2 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[24:23]==2'b11)
      & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_2
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[20:19]==2'b11);
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[22:21]==2'b11);
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_34_2_sdt_1
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[18:17]==2'b11);
  assign c_h_1_5 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_42_4_sdt_4
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[16:15]==2'b11)
      & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_50_2_sdt_2
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[12:11]==2'b11);
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_50_2_sdt_1
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[14:13]==2'b11);
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_58_2_sdt_1
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[10:9]==2'b11);
  assign c_h_1_9 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_50_2_sdt_1
      & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_50_2_sdt_2;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_62_3_sdt_3
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[8:7]==2'b11)
      & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_58_2_sdt_1;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_70_2_sdt_2
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[4:3]==2'b11);
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_70_2_sdt_1
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[6:5]==2'b11);
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_76_2_sdt_1
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[2:1]==2'b11);
  assign c_h_1_12 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_70_2_sdt_1
      & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_42_4_sdt_4;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_90_5_sdt_5
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[0])
      & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_76_2_sdt_1
      & c_h_1_12 & c_h_1_13 & c_h_1_14;
  assign all_same = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_90_5_sdt_5;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_117_nl
      = c_h_1_6 & (c_h_1_13 | (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_42_4_sdt_4));
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_115_nl
      = c_h_1_2 & (c_h_1_5 | (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_62_3_sdt_3))))
      & c_h_1_14));
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_124_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      | (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2))
      & (~((~(out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      & (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_34_2_sdt_1
      | (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_50_2_sdt_1
      & (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_58_2_sdt_1
      | (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_50_2_sdt_2))
      & (~((~(out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_70_2_sdt_1
      & (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_76_2_sdt_1
      | (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14));
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_125_nl
      = (out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[30])
      & ((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[29:28]!=2'b10))
      & (~((~((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[26])
      & ((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[25:24]!=2'b10))))
      & c_h_1_2)) & (~((~((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[22])
      & ((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[21:20]!=2'b10))
      & (~((~((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[18])
      & ((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[17:16]!=2'b10))))
      & c_h_1_5)))) & c_h_1_6)) & (~((~((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[14])
      & ((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[13:12]!=2'b10))
      & (~((~((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[10])
      & ((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[9:8]!=2'b10))))
      & c_h_1_9)) & (~((~((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[6])
      & ((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[5:4]!=2'b10))
      & (~((~((out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_xor_30_0[2:1]==2'b10)))
      & c_h_1_12)))) & c_h_1_13)))) & c_h_1_14));
  assign rtn = MUX_v_5_2_2(({c_h_1_14 , out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_117_nl
      , out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_115_nl ,
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_124_nl , out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_and_125_nl}),
      5'b11111, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_90_5_sdt_5);

  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [30:0] signext_31_1;
    input  vector;
  begin
    signext_31_1= {{30{vector}}, vector};
  end
  endfunction

endmodule




//------> ./GBModule_leading_sign_40_0.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-01
//  Generated date: Wed Feb  4 22:01:35 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_40_0
// ------------------------------------------------------------------


module GBModule_leading_sign_40_0 (
  mantissa, rtn
);
  input [39:0] mantissa;
  output [5:0] rtn;


  // Interconnect Declarations
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_6_2_sdt_2;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_18_3_sdt_3;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_26_2_sdt_2;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_42_4_sdt_4;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_50_2_sdt_2;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_62_3_sdt_3;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_70_2_sdt_2;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_90_5_sdt_5;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_98_2_sdt_2;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_6_2_sdt_1;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_14_2_sdt_1;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_26_2_sdt_1;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_34_2_sdt_1;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_50_2_sdt_1;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_58_2_sdt_1;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_70_2_sdt_1;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_78_2_sdt_1;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_98_2_sdt_1;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_106_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_18;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_155_ssc;

  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_nl;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_or_1_nl;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_2_nl;
  wire[1:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leadi000000;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_nand_nl;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_nand_10_nl;

  // Interconnect Declarations for Component Instantiations
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_6_2_sdt_2
      = ~((mantissa[37:36]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_6_2_sdt_1
      = ~((mantissa[39:38]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_14_2_sdt_1
      = ~((mantissa[35:34]!=2'b00));
  assign c_h_1_2 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_6_2_sdt_1
      & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_6_2_sdt_2;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_18_3_sdt_3
      = (mantissa[33:32]==2'b00) & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_14_2_sdt_1;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_26_2_sdt_2
      = ~((mantissa[29:28]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_26_2_sdt_1
      = ~((mantissa[31:30]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_34_2_sdt_1
      = ~((mantissa[27:26]!=2'b00));
  assign c_h_1_5 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_26_2_sdt_1
      & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_18_3_sdt_3;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_42_4_sdt_4
      = (mantissa[25:24]==2'b00) & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_50_2_sdt_2
      = ~((mantissa[21:20]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_50_2_sdt_1
      = ~((mantissa[23:22]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_58_2_sdt_1
      = ~((mantissa[19:18]!=2'b00));
  assign c_h_1_9 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_50_2_sdt_1
      & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_50_2_sdt_2;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_62_3_sdt_3
      = (mantissa[17:16]==2'b00) & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_58_2_sdt_1;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_70_2_sdt_2
      = ~((mantissa[13:12]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_70_2_sdt_1
      = ~((mantissa[15:14]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_78_2_sdt_1
      = ~((mantissa[11:10]!=2'b00));
  assign c_h_1_12 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_70_2_sdt_1
      & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_42_4_sdt_4;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_90_5_sdt_5
      = (mantissa[9:8]==2'b00) & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_78_2_sdt_1
      & c_h_1_12 & c_h_1_13;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_98_2_sdt_2
      = ~((mantissa[5:4]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_98_2_sdt_1
      = ~((mantissa[7:6]!=2'b00));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_106_2_sdt_1
      = ~((mantissa[3:2]!=2'b00));
  assign c_h_1_17 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_98_2_sdt_1
      & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_98_2_sdt_2;
  assign c_h_1_18 = c_h_1_14 & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_90_5_sdt_5;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_155_ssc
      = (mantissa[1:0]==2'b00) & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_106_2_sdt_1
      & c_h_1_17 & c_h_1_18;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_nl
      = c_h_1_14 & (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_90_5_sdt_5);
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_or_1_nl
      = (c_h_1_6 & (c_h_1_13 | (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_42_4_sdt_4))
      & (~ c_h_1_18)) | ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_155_ssc;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_2_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (c_h_1_17 | (~ c_h_1_18)) & (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_155_ssc);
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_nand_nl
      = ~(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_6_2_sdt_1
      & (ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_14_2_sdt_1
      | (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_26_2_sdt_1
      & (ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_34_2_sdt_1
      | (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_50_2_sdt_1
      & (ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_58_2_sdt_1
      | (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_50_2_sdt_2))
      & (~((~(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_70_2_sdt_1
      & (ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_78_2_sdt_1
      | (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_98_2_sdt_1
      & (ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_106_2_sdt_1
      | (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_wrs_c_98_2_sdt_2))))
      & c_h_1_18)));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_nand_10_nl
      = ~((~((mantissa[39]) | (~((mantissa[38:37]!=2'b01))))) & (~(((mantissa[35])
      | (~((mantissa[34:33]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[31]) | (~((mantissa[30:29]!=2'b01)))))
      & (~(((mantissa[27]) | (~((mantissa[26:25]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[23]) | (~((mantissa[22:21]!=2'b01))))) & (~(((mantissa[19])
      | (~((mantissa[18:17]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[15]) | (~((mantissa[14:13]!=2'b01)))))
      & (~(((mantissa[11]) | (~((mantissa[10:9]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~((~((~((mantissa[7]) | (~((mantissa[6:5]!=2'b01))))) & (~(((mantissa[3])
      | (~((mantissa[2:1]!=2'b01)))) & c_h_1_17)))) & c_h_1_18)));
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leadi000000
      = ~(MUX_v_2_2_2(({ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_nand_nl
      , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_nand_10_nl}),
      2'b11, ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_155_ssc));
  assign rtn = {c_h_1_18 , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_nl
      , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_or_1_nl
      , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_and_2_nl
      , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_leading_1_leadi000000};

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction

endmodule




//------> ./GBModule_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module GBModule_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // spyglass disable SYNTH_5121,W240
    input                s_rst;  // spyglass disable SYNTH_5121,W240
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a; //spyglass disable FlopEConst
                b_reg[0] <= b; //spyglass disable FlopEConst
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> ./GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:55:53 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_is_write_rsc_z, data_memory_index_rsc_z, data_vector_index_rsc_z,
      data_timestep_index_rsc_z, data_write_data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [154:0] this_dat;
  output data_is_write_rsc_z;
  output [1:0] data_memory_index_rsc_z;
  output [7:0] data_vector_index_rsc_z;
  output [15:0] data_timestep_index_rsc_z;
  output [127:0] data_write_data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_data_is_write_rsci_d;
  assign nl_data_is_write_rsci_d = this_dat[0];
  wire [1:0] nl_data_memory_index_rsci_d;
  assign nl_data_memory_index_rsci_d = this_dat[2:1];
  wire [7:0] nl_data_vector_index_rsci_d;
  assign nl_data_vector_index_rsci_d = this_dat[26:19];
  wire [15:0] nl_data_timestep_index_rsci_d;
  assign nl_data_timestep_index_rsci_d = this_dat[18:3];
  wire [127:0] nl_data_write_data_data_rsci_d;
  assign nl_data_write_data_data_rsci_d = this_dat[154:27];
  GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd7),
  .width(32'sd1)) data_is_write_rsci (
      .d(nl_data_is_write_rsci_d),
      .z(data_is_write_rsc_z)
    );
  GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd8),
  .width(32'sd2)) data_memory_index_rsci (
      .d(nl_data_memory_index_rsci_d[1:0]),
      .z(data_memory_index_rsc_z)
    );
  GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd9),
  .width(32'sd8)) data_vector_index_rsci (
      .d(nl_data_vector_index_rsci_d[7:0]),
      .z(data_vector_index_rsc_z)
    );
  GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd10),
  .width(32'sd16)) data_timestep_index_rsci (
      .d(nl_data_timestep_index_rsci_d[15:0]),
      .z(data_timestep_index_rsc_z)
    );
  GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd11),
  .width(32'sd128)) data_write_data_data_rsci (
      .d(nl_data_write_data_data_rsci_d[127:0]),
      .z(data_write_data_data_rsc_z)
    );
  GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd13),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd154),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module GBModule_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_is_write_rsc_z, data_memory_index_rsc_z, data_vector_index_rsc_z,
      data_timestep_index_rsc_z, data_write_data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [154:0] this_dat;
  output data_is_write_rsc_z;
  output [1:0] data_memory_index_rsc_z;
  output [7:0] data_vector_index_rsc_z;
  output [15:0] data_timestep_index_rsc_z;
  output [127:0] data_write_data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_InBlockingless_spec_GB_Large_DataReqcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_is_write_rsc_z(data_is_write_rsc_z),
      .data_memory_index_rsc_z(data_memory_index_rsc_z),
      .data_vector_index_rsc_z(data_vector_index_rsc_z),
      .data_timestep_index_rsc_z(data_timestep_index_rsc_z),
      .data_write_data_data_rsc_z(data_write_data_data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:55:50 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_read_vector_data_data_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [127:0] this_dat;
  reg [127:0] this_dat;
  input [127:0] m_read_vector_data_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [127:0] m_read_vector_data_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd16),
  .width(32'sd128)) m_read_vector_data_data_rsci (
      .dat(m_read_vector_data_data_rsc_dat),
      .idat(m_read_vector_data_data_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd152),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd159)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_read_vector_data_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module GBModule_Connections_OutBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_read_vector_data_data_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [127:0] this_dat;
  input [127:0] m_read_vector_data_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_OutBlockingless_spec_GB_Large_DataRspless_1Ugreater_comma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_read_vector_data_data_rsc_dat(m_read_vector_data_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule_mgc_muladd1_beh.v 
//muladd1
module GBModule_mgc_muladd1(a,b,c,cst,d,z);
  // operation is z = a * (b + d) + c + cst
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_cst = 0;
  parameter signd_cst = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_axb = 1;
  parameter add_c = 1;
  parameter add_d = 1;
  parameter use_const = 1;

  function integer is_square_op;
    input integer alen;
  begin
    if (alen > 1) is_square_op = 0;
    else       is_square_op = 1;
  end endfunction

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_cst-1:0] cst; // spyglass disable SYNTH_5121,W240
  input  [width_d-1:0] d;
  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa;
  reg [width_b-signd_b:0] bb;
  reg [width_c-signd_c:0] cc;
  reg [width_d-signd_d:0] dd;
  reg [width_cst-signd_cst:0] cstin;

  localparam width_bd = (width_d) ? 1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b
                                                                          : width_d - signd_d)
                                  : width_b - signd_b;
  localparam is_square = is_square_op(width_a);
  localparam axb_len = (is_square)?width_bd+1+width_bd+1:width_a-signd_a+1+width_bd+1;

  reg [width_bd:0] bd;
  reg [axb_len-1:0] axb;



  // make all inputs signed
  always @(*) aa = signd_a ? a : {1'b0, a};
  always @(*) bb = signd_b ? b : {1'b0, b};
  generate if (width_c != 0) begin
    always @(*) cc = signd_c ? c : {1'b0, c};
  end endgenerate

  generate if (width_d) begin
    if ( !is_square) begin
      (* keep ="true" *) reg [width_d-signd_d:0] d_keep;
      always @(*) d_keep = signd_d ? d : {1'b0, d};
      always @(*) dd = d_keep;
    end else begin
      always @(*) dd = signd_d ? d : {1'b0, d};
    end
  end endgenerate

  always @(*) cstin = signd_cst ? cst : {1'b0, cst};

  // perform pre-adder
  generate
    if (width_d != 0) begin
      if (add_d) begin always @(*)  bd = $signed(bb) + $signed(dd); end
      else       begin always @(*)  bd = $signed(bb) - $signed(dd); end
    end else     begin always @(*)  bd = $signed(bb); end
  endgenerate

  generate
    if (is_square)
      always @(*) axb = $signed(bd) * $signed(bd);
    else
      always @(*) axb = $signed(aa) * $signed(bd);
  endgenerate

  // perform muladd1
  wire [width_z-1:0]  zz;

  generate
    if (use_const) begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc) + $signed(cstin); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc) + $signed(cstin); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb) + $signed(cstin); end else
      if (!add_axb && !add_c && width_c) begin assign zz = $signed(cstin) - $signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb) + $signed(cstin); end else
                                         begin assign zz = $signed(cstin) - $signed(axb); end
    end  else begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb); end else
      if (!add_axb && !add_c && width_c) begin assign zz = -$signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb); end else
                                         begin assign zz = -$signed(axb); end
    end
  endgenerate

  // adjust output
  assign z = zz;
endmodule // mgc_muladd1

//------> /cad/mentor/2024.2_1/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)
// suppress_sim_read_addr_range_errs:  0 - report errors  1 - suppress errors

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 ,
  parameter suppress_sim_read_addr_range_errs = 1 
  
)( clk,clken,d,q,radr,re,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input  re;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" , syn_ramstyle = "block" *)
  reg [data_width-1:0] mem [depth-1:0];
  integer j;
  initial for (j = 0; j < depth; j = j + 1) mem[j] = 0;
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr READ_ENABLE re
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg re_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
          re_reg <= re;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:55:45 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, m_addr_rsc_dat, m_wstrb_rsc_dat,
      m_rw_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [168:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input [23:0] m_addr_rsc_dat;
  input [15:0] m_wstrb_rsc_dat;
  input m_rw_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [127:0] m_data_rsci_idat;
  wire [23:0] m_addr_rsci_idat;
  wire [15:0] m_wstrb_rsci_idat;
  wire m_rw_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg m_rw_buf_lpi_1_dfm;
  reg [15:0] m_wstrb_buf_lpi_1_dfm;
  reg [23:0] m_addr_buf_lpi_1_dfm;
  reg [127:0] m_data_buf_lpi_1_dfm;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd126),
  .width(32'sd128)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd127),
  .width(32'sd24)) m_addr_rsci (
      .dat(m_addr_rsc_dat),
      .idat(m_addr_rsci_idat)
    );
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd128),
  .width(32'sd16)) m_wstrb_rsci (
      .dat(m_wstrb_rsc_dat),
      .idat(m_wstrb_rsci_idat)
    );
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd129),
  .width(32'sd1)) m_rw_rsci (
      .dat(m_rw_rsc_dat),
      .idat(m_rw_rsci_idat)
    );
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd147),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd156)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = {m_rw_buf_lpi_1_dfm , m_wstrb_buf_lpi_1_dfm , m_addr_buf_lpi_1_dfm
      , m_data_buf_lpi_1_dfm};
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_rw_buf_lpi_1_dfm <= 1'b0;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_rw_buf_lpi_1_dfm <= m_rw_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_wstrb_buf_lpi_1_dfm <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_wstrb_buf_lpi_1_dfm <= m_wstrb_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_addr_buf_lpi_1_dfm <= 24'b000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_addr_buf_lpi_1_dfm <= m_addr_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_lpi_1_dfm <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_lpi_1_dfm <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module GBModule_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, m_addr_rsc_dat, m_wstrb_rsc_dat,
      m_rw_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [168:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input [23:0] m_addr_rsc_dat;
  input [15:0] m_wstrb_rsc_dat;
  input m_rw_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_Push_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_Push_core
      Connections_Combinational_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .m_addr_rsc_dat(m_addr_rsc_dat),
      .m_wstrb_rsc_dat(m_wstrb_rsc_dat),
      .m_rw_rsc_dat(m_rw_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Thu Feb  5 11:55:42 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [127:0] this_dat;
  output [127:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd130),
  .width(32'sd128)) data_data_rsci (
      .d(this_dat),
      .z(data_data_rsc_z)
    );
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd131),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd146),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module GBModule_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [127:0] this_dat;
  output [127:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  GBModule_Connections_Combinationalless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_PopNB_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB_core
      Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./GBModule.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   code@rice-02
//  Generated date: Thu Feb  5 12:25:54 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_RVAOutRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_RVAOutRun_fsm (
  clk, rst, rva_out_Push_mioi_wen_comp, fsm_output
);
  input clk;
  input rst;
  input rva_out_Push_mioi_wen_comp;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for GBModule_GBModule_RVAOutRun_RVAOutRun_fsm_1
  parameter
    RVAOutRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : GBModule_GBModule_RVAOutRun_RVAOutRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // RVAOutRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= RVAOutRun_rlp_C_0;
    end
    else if ( rva_out_Push_mioi_wen_comp ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_staller_1
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_staller_1 (
  clk, rst, RVAOutRun_wten, rva_out_Push_mioi_wen_comp, RVAOutRun_wten_pff
);
  input clk;
  input rst;
  output RVAOutRun_wten;
  input rva_out_Push_mioi_wen_comp;
  output RVAOutRun_wten_pff;


  // Interconnect Declarations
  reg RVAOutRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign RVAOutRun_wten = RVAOutRun_wten_reg;
  assign RVAOutRun_wten_pff = ~ rva_out_Push_mioi_wen_comp;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      RVAOutRun_wten_reg <= 1'b0;
    end
    else begin
      RVAOutRun_wten_reg <= ~ rva_out_Push_mioi_wen_comp;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  RVAOutRun_wen, RVAOutRun_wten, rva_out_Push_mioi_oswt, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_RVAOutRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_oswt_pff
);
  input RVAOutRun_wen;
  input RVAOutRun_wten;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_RVAOutRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & RVAOutRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt)
      & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_RVAOutRun_sct = (~ RVAOutRun_wten)
      & rva_out_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi_nmp_rva_out_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi_nmp_rva_out_PopNB_mio_wait_dp
    (
  clk, rst, nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt, nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt,
      nmp_rva_out_PopNB_mioi_biwt, nmp_rva_out_PopNB_mioi_bdwt, nmp_rva_out_PopNB_mioi_data_data_rsc_z,
      nmp_rva_out_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt;
  output nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt;
  input nmp_rva_out_PopNB_mioi_biwt;
  input nmp_rva_out_PopNB_mioi_bdwt;
  input [127:0] nmp_rva_out_PopNB_mioi_data_data_rsc_z;
  input nmp_rva_out_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg nmp_rva_out_PopNB_mioi_bcwt;
  reg [127:0] nmp_rva_out_PopNB_mioi_data_data_rsc_z_bfwt;
  reg nmp_rva_out_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_128_2_2(nmp_rva_out_PopNB_mioi_data_data_rsc_z,
      nmp_rva_out_PopNB_mioi_data_data_rsc_z_bfwt, nmp_rva_out_PopNB_mioi_bcwt);
  assign nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(nmp_rva_out_PopNB_mioi_return_rsc_z,
      nmp_rva_out_PopNB_mioi_return_rsc_z_bfwt, nmp_rva_out_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_rva_out_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      nmp_rva_out_PopNB_mioi_bcwt <= ~((~(nmp_rva_out_PopNB_mioi_bcwt | nmp_rva_out_PopNB_mioi_biwt))
          | nmp_rva_out_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_rva_out_PopNB_mioi_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      nmp_rva_out_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( nmp_rva_out_PopNB_mioi_biwt ) begin
      nmp_rva_out_PopNB_mioi_data_data_rsc_z_bfwt <= nmp_rva_out_PopNB_mioi_data_data_rsc_z;
      nmp_rva_out_PopNB_mioi_return_rsc_z_bfwt <= nmp_rva_out_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi_nmp_rva_out_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi_nmp_rva_out_PopNB_mio_wait_ctrl
    (
  RVAOutRun_wen, RVAOutRun_wten, nmp_rva_out_PopNB_mioi_oswt, nmp_rva_out_PopNB_mioi_biwt,
      nmp_rva_out_PopNB_mioi_bdwt, nmp_rva_out_PopNB_mioi_biwt_pff, RVAOutRun_wten_pff,
      nmp_rva_out_PopNB_mioi_oswt_pff
);
  input RVAOutRun_wen;
  input RVAOutRun_wten;
  input nmp_rva_out_PopNB_mioi_oswt;
  output nmp_rva_out_PopNB_mioi_biwt;
  output nmp_rva_out_PopNB_mioi_bdwt;
  output nmp_rva_out_PopNB_mioi_biwt_pff;
  input RVAOutRun_wten_pff;
  input nmp_rva_out_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign nmp_rva_out_PopNB_mioi_bdwt = nmp_rva_out_PopNB_mioi_oswt & RVAOutRun_wen;
  assign nmp_rva_out_PopNB_mioi_biwt = (~ RVAOutRun_wten) & nmp_rva_out_PopNB_mioi_oswt;
  assign nmp_rva_out_PopNB_mioi_biwt_pff = (~ RVAOutRun_wten_pff) & nmp_rva_out_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi_gbcore_rva_out_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi_gbcore_rva_out_PopNB_mio_wait_dp
    (
  clk, rst, gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt, gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt,
      gbcore_rva_out_PopNB_mioi_biwt, gbcore_rva_out_PopNB_mioi_bdwt, gbcore_rva_out_PopNB_mioi_data_data_rsc_z,
      gbcore_rva_out_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt;
  output gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt;
  input gbcore_rva_out_PopNB_mioi_biwt;
  input gbcore_rva_out_PopNB_mioi_bdwt;
  input [127:0] gbcore_rva_out_PopNB_mioi_data_data_rsc_z;
  input gbcore_rva_out_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg gbcore_rva_out_PopNB_mioi_bcwt;
  reg [127:0] gbcore_rva_out_PopNB_mioi_data_data_rsc_z_bfwt;
  reg gbcore_rva_out_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_128_2_2(gbcore_rva_out_PopNB_mioi_data_data_rsc_z,
      gbcore_rva_out_PopNB_mioi_data_data_rsc_z_bfwt, gbcore_rva_out_PopNB_mioi_bcwt);
  assign gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(gbcore_rva_out_PopNB_mioi_return_rsc_z,
      gbcore_rva_out_PopNB_mioi_return_rsc_z_bfwt, gbcore_rva_out_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      gbcore_rva_out_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      gbcore_rva_out_PopNB_mioi_bcwt <= ~((~(gbcore_rva_out_PopNB_mioi_bcwt | gbcore_rva_out_PopNB_mioi_biwt))
          | gbcore_rva_out_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      gbcore_rva_out_PopNB_mioi_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      gbcore_rva_out_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( gbcore_rva_out_PopNB_mioi_biwt ) begin
      gbcore_rva_out_PopNB_mioi_data_data_rsc_z_bfwt <= gbcore_rva_out_PopNB_mioi_data_data_rsc_z;
      gbcore_rva_out_PopNB_mioi_return_rsc_z_bfwt <= gbcore_rva_out_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi_gbcore_rva_out_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi_gbcore_rva_out_PopNB_mio_wait_ctrl
    (
  RVAOutRun_wen, RVAOutRun_wten, gbcore_rva_out_PopNB_mioi_oswt, gbcore_rva_out_PopNB_mioi_biwt,
      gbcore_rva_out_PopNB_mioi_bdwt, gbcore_rva_out_PopNB_mioi_biwt_pff, RVAOutRun_wten_pff,
      gbcore_rva_out_PopNB_mioi_oswt_pff
);
  input RVAOutRun_wen;
  input RVAOutRun_wten;
  input gbcore_rva_out_PopNB_mioi_oswt;
  output gbcore_rva_out_PopNB_mioi_biwt;
  output gbcore_rva_out_PopNB_mioi_bdwt;
  output gbcore_rva_out_PopNB_mioi_biwt_pff;
  input RVAOutRun_wten_pff;
  input gbcore_rva_out_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign gbcore_rva_out_PopNB_mioi_bdwt = gbcore_rva_out_PopNB_mioi_oswt & RVAOutRun_wen;
  assign gbcore_rva_out_PopNB_mioi_biwt = (~ RVAOutRun_wten) & gbcore_rva_out_PopNB_mioi_oswt;
  assign gbcore_rva_out_PopNB_mioi_biwt_pff = (~ RVAOutRun_wten_pff) & gbcore_rva_out_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_RVAInRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_RVAInRun_fsm (
  clk, rst, RVAInRun_wen, fsm_output
);
  input clk;
  input rst;
  input RVAInRun_wen;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for GBModule_GBModule_RVAInRun_RVAInRun_fsm_1
  parameter
    RVAInRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : GBModule_GBModule_RVAInRun_RVAInRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // RVAInRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= RVAInRun_rlp_C_0;
    end
    else if ( RVAInRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_staller
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_staller (
  clk, rst, RVAInRun_wen, RVAInRun_wten, gbcore_rva_in_Push_mioi_wen_comp, nmp_rva_in_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output RVAInRun_wen;
  output RVAInRun_wten;
  input gbcore_rva_in_Push_mioi_wen_comp;
  input nmp_rva_in_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg RVAInRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign RVAInRun_wen = gbcore_rva_in_Push_mioi_wen_comp & nmp_rva_in_Push_mioi_wen_comp;
  assign RVAInRun_wten = RVAInRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      RVAInRun_wten_reg <= 1'b0;
    end
    else begin
      RVAInRun_wten_reg <= ~ RVAInRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_dp
    (
  clk, rst, nmp_rva_in_Push_mioi_oswt, nmp_rva_in_Push_mioi_wen_comp, nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun,
      nmp_rva_in_Push_mioi_biwt, nmp_rva_in_Push_mioi_bdwt, nmp_rva_in_Push_mioi_bcwt,
      nmp_rva_in_Push_mioi_m_addr_rsc_dat
);
  input clk;
  input rst;
  input nmp_rva_in_Push_mioi_oswt;
  output nmp_rva_in_Push_mioi_wen_comp;
  input [23:0] nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun;
  input nmp_rva_in_Push_mioi_biwt;
  input nmp_rva_in_Push_mioi_bdwt;
  output nmp_rva_in_Push_mioi_bcwt;
  reg nmp_rva_in_Push_mioi_bcwt;
  output [23:0] nmp_rva_in_Push_mioi_m_addr_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  assign nmp_rva_in_Push_mioi_wen_comp = (~ nmp_rva_in_Push_mioi_oswt) | nmp_rva_in_Push_mioi_biwt
      | nmp_rva_in_Push_mioi_bcwt;
  assign nmp_rva_in_Push_mioi_m_addr_rsc_dat = {4'b1100 , (nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun[19:0])};
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_rva_in_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      nmp_rva_in_Push_mioi_bcwt <= ~((~(nmp_rva_in_Push_mioi_bcwt | nmp_rva_in_Push_mioi_biwt))
          | nmp_rva_in_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_ctrl
    (
  RVAInRun_wen, nmp_rva_in_Push_mioi_oswt, nmp_rva_in_Push_mioi_biwt, nmp_rva_in_Push_mioi_bdwt,
      nmp_rva_in_Push_mioi_bcwt, nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct,
      nmp_rva_in_Push_mioi_ccs_ccore_done_sync_vld, nmp_rva_in_Push_mioi_oswt_pff
);
  input RVAInRun_wen;
  input nmp_rva_in_Push_mioi_oswt;
  output nmp_rva_in_Push_mioi_biwt;
  output nmp_rva_in_Push_mioi_bdwt;
  input nmp_rva_in_Push_mioi_bcwt;
  output nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct;
  input nmp_rva_in_Push_mioi_ccs_ccore_done_sync_vld;
  input nmp_rva_in_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign nmp_rva_in_Push_mioi_bdwt = nmp_rva_in_Push_mioi_oswt & RVAInRun_wen;
  assign nmp_rva_in_Push_mioi_biwt = nmp_rva_in_Push_mioi_oswt & (~ nmp_rva_in_Push_mioi_bcwt)
      & nmp_rva_in_Push_mioi_ccs_ccore_done_sync_vld;
  assign nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct = RVAInRun_wen & nmp_rva_in_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_gbcore_rva_in_Push_mioi_gbcore_rva_in_Push_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_gbcore_rva_in_Push_mioi_gbcore_rva_in_Push_mio_wait_dp
    (
  clk, rst, gbcore_rva_in_Push_mioi_oswt, gbcore_rva_in_Push_mioi_wen_comp, gbcore_rva_in_Push_mioi_biwt,
      gbcore_rva_in_Push_mioi_bdwt, gbcore_rva_in_Push_mioi_bcwt
);
  input clk;
  input rst;
  input gbcore_rva_in_Push_mioi_oswt;
  output gbcore_rva_in_Push_mioi_wen_comp;
  input gbcore_rva_in_Push_mioi_biwt;
  input gbcore_rva_in_Push_mioi_bdwt;
  output gbcore_rva_in_Push_mioi_bcwt;
  reg gbcore_rva_in_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign gbcore_rva_in_Push_mioi_wen_comp = (~ gbcore_rva_in_Push_mioi_oswt) | gbcore_rva_in_Push_mioi_biwt
      | gbcore_rva_in_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      gbcore_rva_in_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      gbcore_rva_in_Push_mioi_bcwt <= ~((~(gbcore_rva_in_Push_mioi_bcwt | gbcore_rva_in_Push_mioi_biwt))
          | gbcore_rva_in_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_gbcore_rva_in_Push_mioi_gbcore_rva_in_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_gbcore_rva_in_Push_mioi_gbcore_rva_in_Push_mio_wait_ctrl
    (
  RVAInRun_wen, gbcore_rva_in_Push_mioi_oswt, gbcore_rva_in_Push_mioi_biwt, gbcore_rva_in_Push_mioi_bdwt,
      gbcore_rva_in_Push_mioi_bcwt, gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct,
      gbcore_rva_in_Push_mioi_ccs_ccore_done_sync_vld, gbcore_rva_in_Push_mioi_oswt_pff
);
  input RVAInRun_wen;
  input gbcore_rva_in_Push_mioi_oswt;
  output gbcore_rva_in_Push_mioi_biwt;
  output gbcore_rva_in_Push_mioi_bdwt;
  input gbcore_rva_in_Push_mioi_bcwt;
  output gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct;
  input gbcore_rva_in_Push_mioi_ccs_ccore_done_sync_vld;
  input gbcore_rva_in_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign gbcore_rva_in_Push_mioi_bdwt = gbcore_rva_in_Push_mioi_oswt & RVAInRun_wen;
  assign gbcore_rva_in_Push_mioi_biwt = gbcore_rva_in_Push_mioi_oswt & (~ gbcore_rva_in_Push_mioi_bcwt)
      & gbcore_rva_in_Push_mioi_ccs_ccore_done_sync_vld;
  assign gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct = RVAInRun_wen & gbcore_rva_in_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt,
      rva_in_PopNB_mioi_return_rsc_z_mxwt, rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt,
      rva_in_PopNB_mioi_data_data_rsc_z, rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_wstrb_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [23:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output [15:0] rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input [15:0] rva_in_PopNB_mioi_data_wstrb_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [127:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg [23:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt;
  reg [15:0] rva_in_PopNB_mioi_data_wstrb_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_128_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_24_2_2(rva_in_PopNB_mioi_data_addr_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt = MUX_v_16_2_2(rva_in_PopNB_mioi_data_wstrb_rsc_z,
      rva_in_PopNB_mioi_data_wstrb_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt <= 24'b000000000000000000000000;
      rva_in_PopNB_mioi_data_wstrb_rsc_z_bfwt <= 16'b0000000000000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt <= rva_in_PopNB_mioi_data_addr_rsc_z;
      rva_in_PopNB_mioi_data_wstrb_rsc_z_bfwt <= rva_in_PopNB_mioi_data_wstrb_rsc_z;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [23:0] MUX_v_24_2_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input  sel;
    reg [23:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_24_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  RVAInRun_wen, RVAInRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt,
      rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input RVAInRun_wen;
  input RVAInRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & RVAInRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ RVAInRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = RVAInRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_77_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_77_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_76_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_76_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_75_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_75_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_74_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_74_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_73_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_73_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_72_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_72_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_71_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_71_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_70_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_70_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_69_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_69_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_68_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_68_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_67_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_67_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_66_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_66_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_65_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_65_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_64_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_64_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_63_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_63_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_62_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_62_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_GBCoreRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_GBCoreRun_fsm (
  clk, rst, GBCoreRun_wen, fsm_output
);
  input clk;
  input rst;
  input GBCoreRun_wen;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for GBModule_GBCore_GBCoreRun_GBCoreRun_fsm_1
  parameter
    GBCoreRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : GBModule_GBCore_GBCoreRun_GBCoreRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // GBCoreRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= GBCoreRun_rlp_C_0;
    end
    else if ( GBCoreRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_staller
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_staller (
  clk, rst, GBCoreRun_wen, GBCoreRun_wten, rva_out_large_Push_mioi_wen_comp, nmp_large_rsp_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output GBCoreRun_wen;
  output GBCoreRun_wten;
  input rva_out_large_Push_mioi_wen_comp;
  input nmp_large_rsp_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg GBCoreRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign GBCoreRun_wen = rva_out_large_Push_mioi_wen_comp & nmp_large_rsp_Push_mioi_wen_comp;
  assign GBCoreRun_wten = GBCoreRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCoreRun_wten_reg <= 1'b0;
    end
    else begin
      GBCoreRun_wten_reg <= ~ GBCoreRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_wait_dp
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_wait_dp (
  large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d, large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d,
      large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d, large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d,
      large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d, large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d,
      large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d, large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d,
      large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d, large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d,
      large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d, large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d,
      large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d, large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d,
      large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d, large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d,
      GBCoreRun_wen, large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo, large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo, large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo, large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo, large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo, large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo, large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo, large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo, large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo, large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo, large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo, large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo, large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo, large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo, large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo, large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo_ir_unreg,
      large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo, large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo_ir_unreg
);
  output large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d;
  output large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d;
  output large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d;
  output large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d;
  output large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d;
  output large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d;
  output large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d;
  output large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d;
  output large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d;
  output large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d;
  output large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d;
  output large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d;
  output large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d;
  output large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d;
  output large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d;
  output large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d;
  input GBCoreRun_wen;
  input large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo;
  input large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo;
  input large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo;
  input large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo;
  input large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo;
  input large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo;
  input large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo;
  input large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo;
  input large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo;
  input large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo;
  input large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo;
  input large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo;
  input large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo;
  input large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo;
  input large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo;
  input large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo_ir_unreg;
  input large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo;
  input large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo_ir_unreg;



  // Interconnect Declarations for Component Instantiations 
  assign large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo
      | large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo
      | large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo
      | large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo
      | large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo
      | large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo
      | large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo
      | large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo
      | large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo
      | large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo
      | large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo
      | large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo
      | large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo
      | large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo
      | large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo
      | large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo_ir_unreg);
  assign large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d = GBCoreRun_wen & (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo
      | large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo_ir_unreg);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_nmp_large_rsp_Push_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_nmp_large_rsp_Push_mio_wait_dp
    (
  clk, rst, nmp_large_rsp_Push_mioi_oswt, nmp_large_rsp_Push_mioi_wen_comp, nmp_large_rsp_Push_mioi_biwt,
      nmp_large_rsp_Push_mioi_bdwt, nmp_large_rsp_Push_mioi_bcwt
);
  input clk;
  input rst;
  input nmp_large_rsp_Push_mioi_oswt;
  output nmp_large_rsp_Push_mioi_wen_comp;
  input nmp_large_rsp_Push_mioi_biwt;
  input nmp_large_rsp_Push_mioi_bdwt;
  output nmp_large_rsp_Push_mioi_bcwt;
  reg nmp_large_rsp_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign nmp_large_rsp_Push_mioi_wen_comp = (~ nmp_large_rsp_Push_mioi_oswt) | nmp_large_rsp_Push_mioi_biwt
      | nmp_large_rsp_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_large_rsp_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      nmp_large_rsp_Push_mioi_bcwt <= ~((~(nmp_large_rsp_Push_mioi_bcwt | nmp_large_rsp_Push_mioi_biwt))
          | nmp_large_rsp_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_nmp_large_rsp_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_nmp_large_rsp_Push_mio_wait_ctrl
    (
  GBCoreRun_wen, nmp_large_rsp_Push_mioi_oswt, nmp_large_rsp_Push_mioi_biwt, nmp_large_rsp_Push_mioi_bdwt,
      nmp_large_rsp_Push_mioi_bcwt, nmp_large_rsp_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct,
      nmp_large_rsp_Push_mioi_ccs_ccore_done_sync_vld, nmp_large_rsp_Push_mioi_oswt_pff
);
  input GBCoreRun_wen;
  input nmp_large_rsp_Push_mioi_oswt;
  output nmp_large_rsp_Push_mioi_biwt;
  output nmp_large_rsp_Push_mioi_bdwt;
  input nmp_large_rsp_Push_mioi_bcwt;
  output nmp_large_rsp_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct;
  input nmp_large_rsp_Push_mioi_ccs_ccore_done_sync_vld;
  input nmp_large_rsp_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign nmp_large_rsp_Push_mioi_bdwt = nmp_large_rsp_Push_mioi_oswt & GBCoreRun_wen;
  assign nmp_large_rsp_Push_mioi_biwt = nmp_large_rsp_Push_mioi_oswt & (~ nmp_large_rsp_Push_mioi_bcwt)
      & nmp_large_rsp_Push_mioi_ccs_ccore_done_sync_vld;
  assign nmp_large_rsp_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct = GBCoreRun_wen
      & nmp_large_rsp_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_rva_out_large_Push_mioi_rva_out_large_Push_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_rva_out_large_Push_mioi_rva_out_large_Push_mio_wait_dp
    (
  clk, rst, rva_out_large_Push_mioi_oswt, rva_out_large_Push_mioi_wen_comp, rva_out_large_Push_mioi_biwt,
      rva_out_large_Push_mioi_bdwt, rva_out_large_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_large_Push_mioi_oswt;
  output rva_out_large_Push_mioi_wen_comp;
  input rva_out_large_Push_mioi_biwt;
  input rva_out_large_Push_mioi_bdwt;
  output rva_out_large_Push_mioi_bcwt;
  reg rva_out_large_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_large_Push_mioi_wen_comp = (~ rva_out_large_Push_mioi_oswt) | rva_out_large_Push_mioi_biwt
      | rva_out_large_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_large_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_large_Push_mioi_bcwt <= ~((~(rva_out_large_Push_mioi_bcwt | rva_out_large_Push_mioi_biwt))
          | rva_out_large_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_rva_out_large_Push_mioi_rva_out_large_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_rva_out_large_Push_mioi_rva_out_large_Push_mio_wait_ctrl
    (
  GBCoreRun_wen, rva_out_large_Push_mioi_oswt, rva_out_large_Push_mioi_biwt, rva_out_large_Push_mioi_bdwt,
      rva_out_large_Push_mioi_bcwt, rva_out_large_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct,
      rva_out_large_Push_mioi_ccs_ccore_done_sync_vld, rva_out_large_Push_mioi_oswt_pff
);
  input GBCoreRun_wen;
  input rva_out_large_Push_mioi_oswt;
  output rva_out_large_Push_mioi_biwt;
  output rva_out_large_Push_mioi_bdwt;
  input rva_out_large_Push_mioi_bcwt;
  output rva_out_large_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct;
  input rva_out_large_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_large_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_large_Push_mioi_bdwt = rva_out_large_Push_mioi_oswt & GBCoreRun_wen;
  assign rva_out_large_Push_mioi_biwt = rva_out_large_Push_mioi_oswt & (~ rva_out_large_Push_mioi_bcwt)
      & rva_out_large_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_large_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct = GBCoreRun_wen
      & rva_out_large_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_nmp_large_req_PopNB_mioi_nmp_large_req_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_nmp_large_req_PopNB_mioi_nmp_large_req_PopNB_mio_wait_dp
    (
  clk, rst, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt, nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt,
      nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt, nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt,
      nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt,
      nmp_large_req_PopNB_mioi_biwt, nmp_large_req_PopNB_mioi_bdwt, nmp_large_req_PopNB_mioi_data_is_write_rsc_z,
      nmp_large_req_PopNB_mioi_data_memory_index_rsc_z, nmp_large_req_PopNB_mioi_data_vector_index_rsc_z,
      nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z, nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z,
      nmp_large_req_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt;
  output [1:0] nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt;
  output [7:0] nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt;
  output [15:0] nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt;
  output [127:0] nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt;
  output nmp_large_req_PopNB_mioi_return_rsc_z_mxwt;
  input nmp_large_req_PopNB_mioi_biwt;
  input nmp_large_req_PopNB_mioi_bdwt;
  input nmp_large_req_PopNB_mioi_data_is_write_rsc_z;
  input [1:0] nmp_large_req_PopNB_mioi_data_memory_index_rsc_z;
  input [7:0] nmp_large_req_PopNB_mioi_data_vector_index_rsc_z;
  input [15:0] nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z;
  input [127:0] nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z;
  input nmp_large_req_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg nmp_large_req_PopNB_mioi_bcwt;
  reg nmp_large_req_PopNB_mioi_data_is_write_rsc_z_bfwt;
  reg [1:0] nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_bfwt;
  reg [7:0] nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_bfwt;
  reg [15:0] nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_bfwt;
  reg [127:0] nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_bfwt;
  reg nmp_large_req_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt = MUX_s_1_2_2(nmp_large_req_PopNB_mioi_data_is_write_rsc_z,
      nmp_large_req_PopNB_mioi_data_is_write_rsc_z_bfwt, nmp_large_req_PopNB_mioi_bcwt);
  assign nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt = MUX_v_2_2_2(nmp_large_req_PopNB_mioi_data_memory_index_rsc_z,
      nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_bfwt, nmp_large_req_PopNB_mioi_bcwt);
  assign nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt = MUX_v_8_2_2(nmp_large_req_PopNB_mioi_data_vector_index_rsc_z,
      nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_bfwt, nmp_large_req_PopNB_mioi_bcwt);
  assign nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt = MUX_v_16_2_2(nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z,
      nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_bfwt, nmp_large_req_PopNB_mioi_bcwt);
  assign nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt = MUX_v_128_2_2(nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z,
      nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_bfwt, nmp_large_req_PopNB_mioi_bcwt);
  assign nmp_large_req_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(nmp_large_req_PopNB_mioi_return_rsc_z,
      nmp_large_req_PopNB_mioi_return_rsc_z_bfwt, nmp_large_req_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_large_req_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      nmp_large_req_PopNB_mioi_bcwt <= ~((~(nmp_large_req_PopNB_mioi_bcwt | nmp_large_req_PopNB_mioi_biwt))
          | nmp_large_req_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_large_req_PopNB_mioi_data_is_write_rsc_z_bfwt <= 1'b0;
      nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_bfwt <= 2'b00;
      nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_bfwt <= 8'b00000000;
      nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_bfwt <= 16'b0000000000000000;
      nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      nmp_large_req_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( nmp_large_req_PopNB_mioi_biwt ) begin
      nmp_large_req_PopNB_mioi_data_is_write_rsc_z_bfwt <= nmp_large_req_PopNB_mioi_data_is_write_rsc_z;
      nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_bfwt <= nmp_large_req_PopNB_mioi_data_memory_index_rsc_z;
      nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_bfwt <= nmp_large_req_PopNB_mioi_data_vector_index_rsc_z;
      nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_bfwt <= nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z;
      nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_bfwt <= nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z;
      nmp_large_req_PopNB_mioi_return_rsc_z_bfwt <= nmp_large_req_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_nmp_large_req_PopNB_mioi_nmp_large_req_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_nmp_large_req_PopNB_mioi_nmp_large_req_PopNB_mio_wait_ctrl
    (
  GBCoreRun_wen, GBCoreRun_wten, nmp_large_req_PopNB_mioi_oswt, nmp_large_req_PopNB_mioi_biwt,
      nmp_large_req_PopNB_mioi_bdwt, nmp_large_req_PopNB_mioi_biwt_pff, nmp_large_req_PopNB_mioi_oswt_pff
);
  input GBCoreRun_wen;
  input GBCoreRun_wten;
  input nmp_large_req_PopNB_mioi_oswt;
  output nmp_large_req_PopNB_mioi_biwt;
  output nmp_large_req_PopNB_mioi_bdwt;
  output nmp_large_req_PopNB_mioi_biwt_pff;
  input nmp_large_req_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign nmp_large_req_PopNB_mioi_bdwt = nmp_large_req_PopNB_mioi_oswt & GBCoreRun_wen;
  assign nmp_large_req_PopNB_mioi_biwt = (~ GBCoreRun_wten) & nmp_large_req_PopNB_mioi_oswt;
  assign nmp_large_req_PopNB_mioi_biwt_pff = GBCoreRun_wen & nmp_large_req_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_rva_in_large_PopNB_mioi_rva_in_large_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_rva_in_large_PopNB_mioi_rva_in_large_PopNB_mio_wait_dp
    (
  clk, rst, rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_large_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_large_PopNB_mioi_biwt, rva_in_large_PopNB_mioi_bdwt, rva_in_large_PopNB_mioi_data_data_rsc_z,
      rva_in_large_PopNB_mioi_data_addr_rsc_z, rva_in_large_PopNB_mioi_data_rw_rsc_z,
      rva_in_large_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_large_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_large_PopNB_mioi_biwt;
  input rva_in_large_PopNB_mioi_bdwt;
  input [127:0] rva_in_large_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_large_PopNB_mioi_data_addr_rsc_z;
  input rva_in_large_PopNB_mioi_data_rw_rsc_z;
  input rva_in_large_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_large_PopNB_mioi_bcwt;
  reg [127:0] rva_in_large_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_large_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_large_PopNB_mioi_return_rsc_z_bfwt;
  reg [19:0] rva_in_large_PopNB_mioi_data_addr_rsc_z_bfwt_23_4;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_128_2_2(rva_in_large_PopNB_mioi_data_data_rsc_z,
      rva_in_large_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_large_PopNB_mioi_bcwt);
  assign rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_large_PopNB_mioi_data_rw_rsc_z,
      rva_in_large_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_large_PopNB_mioi_bcwt);
  assign rva_in_large_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_large_PopNB_mioi_return_rsc_z,
      rva_in_large_PopNB_mioi_return_rsc_z_bfwt, rva_in_large_PopNB_mioi_bcwt);
  assign rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_20_2_2((rva_in_large_PopNB_mioi_data_addr_rsc_z[23:4]),
      rva_in_large_PopNB_mioi_data_addr_rsc_z_bfwt_23_4, rva_in_large_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_large_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_large_PopNB_mioi_bcwt <= ~((~(rva_in_large_PopNB_mioi_bcwt | rva_in_large_PopNB_mioi_biwt))
          | rva_in_large_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_large_PopNB_mioi_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_large_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= 20'b00000000000000000000;
      rva_in_large_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_large_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_large_PopNB_mioi_biwt ) begin
      rva_in_large_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_large_PopNB_mioi_data_data_rsc_z;
      rva_in_large_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= rva_in_large_PopNB_mioi_data_addr_rsc_z[23:4];
      rva_in_large_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_large_PopNB_mioi_data_rw_rsc_z;
      rva_in_large_PopNB_mioi_return_rsc_z_bfwt <= rva_in_large_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_rva_in_large_PopNB_mioi_rva_in_large_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_rva_in_large_PopNB_mioi_rva_in_large_PopNB_mio_wait_ctrl
    (
  GBCoreRun_wen, GBCoreRun_wten, rva_in_large_PopNB_mioi_oswt, rva_in_large_PopNB_mioi_biwt,
      rva_in_large_PopNB_mioi_bdwt, rva_in_large_PopNB_mioi_biwt_pff, rva_in_large_PopNB_mioi_oswt_pff
);
  input GBCoreRun_wen;
  input GBCoreRun_wten;
  input rva_in_large_PopNB_mioi_oswt;
  output rva_in_large_PopNB_mioi_biwt;
  output rva_in_large_PopNB_mioi_bdwt;
  output rva_in_large_PopNB_mioi_biwt_pff;
  input rva_in_large_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_large_PopNB_mioi_bdwt = rva_in_large_PopNB_mioi_oswt & GBCoreRun_wen;
  assign rva_in_large_PopNB_mioi_biwt = (~ GBCoreRun_wten) & rva_in_large_PopNB_mioi_oswt;
  assign rva_in_large_PopNB_mioi_biwt_pff = GBCoreRun_wen & rva_in_large_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_NMPRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_NMPRun_fsm (
  clk, rst, NMPRun_wen, fsm_output
);
  input clk;
  input rst;
  input NMPRun_wen;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for GBModule_NMP_NMPRun_NMPRun_fsm_1
  parameter
    NMPRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : GBModule_NMP_NMPRun_NMPRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // NMPRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= NMPRun_rlp_C_0;
    end
    else if ( NMPRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_staller
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_staller (
  clk, rst, NMPRun_wen, NMPRun_wten, large_req_Push_mioi_wen_comp, rva_out_Push_mioi_wen_comp,
      done_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output NMPRun_wen;
  output NMPRun_wten;
  input large_req_Push_mioi_wen_comp;
  input rva_out_Push_mioi_wen_comp;
  input done_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg NMPRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign NMPRun_wen = large_req_Push_mioi_wen_comp & rva_out_Push_mioi_wen_comp &
      done_Push_mioi_wen_comp;
  assign NMPRun_wten = NMPRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMPRun_wten_reg <= 1'b0;
    end
    else begin
      NMPRun_wten_reg <= ~ NMPRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_wait_dp
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_wait_dp (
  NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_en, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en,
      NMPRun_wen, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo_ir_unreg,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo_ir_unreg,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo, NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo_ir_unreg,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo_ir_unreg
);
  output NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en;
  output NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en;
  output NMP_ComputeRMSNormalize_for_1_mul_cmp_en;
  output NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en;
  input NMPRun_wen;
  input NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo;
  input NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo_ir_unreg;
  input NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo;
  input NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo_ir_unreg;
  input NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo;
  input NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo_ir_unreg;
  input NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo;
  input NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo_ir_unreg;



  // Interconnect Declarations for Component Instantiations 
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en = NMPRun_wen & (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo
      | NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo_ir_unreg);
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en
      = NMPRun_wen & (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo
      | NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo_ir_unreg);
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_en = NMPRun_wen & (NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo
      | NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo_ir_unreg);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en = NMPRun_wen
      & (NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo | NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo_ir_unreg);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_done_Push_mioi_done_Push_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_done_Push_mioi_done_Push_mio_wait_dp (
  clk, rst, done_Push_mioi_oswt, done_Push_mioi_wen_comp, done_Push_mioi_biwt, done_Push_mioi_bdwt,
      done_Push_mioi_bcwt
);
  input clk;
  input rst;
  input done_Push_mioi_oswt;
  output done_Push_mioi_wen_comp;
  input done_Push_mioi_biwt;
  input done_Push_mioi_bdwt;
  output done_Push_mioi_bcwt;
  reg done_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_Push_mioi_wen_comp = (~ done_Push_mioi_oswt) | done_Push_mioi_biwt
      | done_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      done_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      done_Push_mioi_bcwt <= ~((~(done_Push_mioi_bcwt | done_Push_mioi_biwt)) | done_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_done_Push_mioi_done_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_done_Push_mioi_done_Push_mio_wait_ctrl (
  NMPRun_wen, done_Push_mioi_oswt, done_Push_mioi_biwt, done_Push_mioi_bdwt, done_Push_mioi_bcwt,
      done_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct, done_Push_mioi_ccs_ccore_done_sync_vld,
      done_Push_mioi_oswt_pff
);
  input NMPRun_wen;
  input done_Push_mioi_oswt;
  output done_Push_mioi_biwt;
  output done_Push_mioi_bdwt;
  input done_Push_mioi_bcwt;
  output done_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct;
  input done_Push_mioi_ccs_ccore_done_sync_vld;
  input done_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign done_Push_mioi_bdwt = done_Push_mioi_oswt & NMPRun_wen;
  assign done_Push_mioi_biwt = done_Push_mioi_oswt & (~ done_Push_mioi_bcwt) & done_Push_mioi_ccs_ccore_done_sync_vld;
  assign done_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct = NMPRun_wen & done_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt, rva_out_Push_mioi_m_data_rsc_dat,
      rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;
  output [127:0] rva_out_Push_mioi_m_data_rsc_dat;
  input [127:0] rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  assign rva_out_Push_mioi_m_data_rsc_dat = {29'b00000000000000000000000000000 ,
      (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[98:96]) , 16'b0000000000000000
      , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[79:64]) , 8'b00000000 , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[55:48])
      , 13'b0000000000000 , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[34:32])
      , 21'b000000000000000000000 , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[10:8])
      , 7'b0000000 , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[0])};
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  NMPRun_wen, rva_out_Push_mioi_oswt, rva_out_Push_mioi_biwt, rva_out_Push_mioi_bdwt,
      rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_oswt_pff
);
  input NMPRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & NMPRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt)
      & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct = NMPRun_wen & rva_out_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_large_rsp_PopNB_mioi_large_rsp_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_large_rsp_PopNB_mioi_large_rsp_PopNB_mio_wait_dp (
  clk, rst, large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt, large_rsp_PopNB_mioi_return_rsc_z_mxwt,
      large_rsp_PopNB_mioi_biwt, large_rsp_PopNB_mioi_bdwt, large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z,
      large_rsp_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt;
  output large_rsp_PopNB_mioi_return_rsc_z_mxwt;
  input large_rsp_PopNB_mioi_biwt;
  input large_rsp_PopNB_mioi_bdwt;
  input [127:0] large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z;
  input large_rsp_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg large_rsp_PopNB_mioi_bcwt;
  reg [127:0] large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_bfwt;
  reg large_rsp_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt = MUX_v_128_2_2(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z,
      large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_bfwt, large_rsp_PopNB_mioi_bcwt);
  assign large_rsp_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(large_rsp_PopNB_mioi_return_rsc_z,
      large_rsp_PopNB_mioi_return_rsc_z_bfwt, large_rsp_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_rsp_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      large_rsp_PopNB_mioi_bcwt <= ~((~(large_rsp_PopNB_mioi_bcwt | large_rsp_PopNB_mioi_biwt))
          | large_rsp_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      large_rsp_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( large_rsp_PopNB_mioi_biwt ) begin
      large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_bfwt <= large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z;
      large_rsp_PopNB_mioi_return_rsc_z_bfwt <= large_rsp_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_large_rsp_PopNB_mioi_large_rsp_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_large_rsp_PopNB_mioi_large_rsp_PopNB_mio_wait_ctrl (
  NMPRun_wen, NMPRun_wten, large_rsp_PopNB_mioi_oswt, large_rsp_PopNB_mioi_biwt,
      large_rsp_PopNB_mioi_bdwt, large_rsp_PopNB_mioi_biwt_pff, large_rsp_PopNB_mioi_oswt_pff
);
  input NMPRun_wen;
  input NMPRun_wten;
  input large_rsp_PopNB_mioi_oswt;
  output large_rsp_PopNB_mioi_biwt;
  output large_rsp_PopNB_mioi_bdwt;
  output large_rsp_PopNB_mioi_biwt_pff;
  input large_rsp_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign large_rsp_PopNB_mioi_bdwt = large_rsp_PopNB_mioi_oswt & NMPRun_wen;
  assign large_rsp_PopNB_mioi_biwt = (~ NMPRun_wten) & large_rsp_PopNB_mioi_oswt;
  assign large_rsp_PopNB_mioi_biwt_pff = NMPRun_wen & large_rsp_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  NMPRun_wen, NMPRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt,
      start_PopNB_mioi_biwt_pff, start_PopNB_mioi_oswt_pff
);
  input NMPRun_wen;
  input NMPRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_biwt_pff;
  input start_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & NMPRun_wen;
  assign start_PopNB_mioi_biwt = (~ NMPRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_biwt_pff = NMPRun_wen & start_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_large_req_Push_mioi_large_req_Push_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_large_req_Push_mioi_large_req_Push_mio_wait_dp (
  clk, rst, large_req_Push_mioi_oswt, large_req_Push_mioi_wen_comp, large_req_Push_mioi_biwt,
      large_req_Push_mioi_bdwt, large_req_Push_mioi_bcwt
);
  input clk;
  input rst;
  input large_req_Push_mioi_oswt;
  output large_req_Push_mioi_wen_comp;
  input large_req_Push_mioi_biwt;
  input large_req_Push_mioi_bdwt;
  output large_req_Push_mioi_bcwt;
  reg large_req_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign large_req_Push_mioi_wen_comp = (~ large_req_Push_mioi_oswt) | large_req_Push_mioi_biwt
      | large_req_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_req_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      large_req_Push_mioi_bcwt <= ~((~(large_req_Push_mioi_bcwt | large_req_Push_mioi_biwt))
          | large_req_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_large_req_Push_mioi_large_req_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_large_req_Push_mioi_large_req_Push_mio_wait_ctrl (
  NMPRun_wen, large_req_Push_mioi_oswt, large_req_Push_mioi_biwt, large_req_Push_mioi_bdwt,
      large_req_Push_mioi_bcwt, large_req_Push_mioi_m_is_write_rsc_dat_NMPRun_sct,
      large_req_Push_mioi_ccs_ccore_done_sync_vld, large_req_Push_mioi_oswt_pff
);
  input NMPRun_wen;
  input large_req_Push_mioi_oswt;
  output large_req_Push_mioi_biwt;
  output large_req_Push_mioi_bdwt;
  input large_req_Push_mioi_bcwt;
  output large_req_Push_mioi_m_is_write_rsc_dat_NMPRun_sct;
  input large_req_Push_mioi_ccs_ccore_done_sync_vld;
  input large_req_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign large_req_Push_mioi_bdwt = large_req_Push_mioi_oswt & NMPRun_wen;
  assign large_req_Push_mioi_biwt = large_req_Push_mioi_oswt & (~ large_req_Push_mioi_bcwt)
      & large_req_Push_mioi_ccs_ccore_done_sync_vld;
  assign large_req_Push_mioi_m_is_write_rsc_dat_NMPRun_sct = NMPRun_wen & large_req_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [33:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  reg [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4;
  reg [2:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt_98_96;
  reg [15:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt_79_64;
  reg [7:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt_55_48;
  reg [2:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt_34_32;
  reg [2:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt_10_8;
  reg rva_in_PopNB_mioi_data_data_rsc_z_bfwt_0;

  wire[2:0] while_if_mux_1_nl;
  wire[15:0] while_if_mux_11_nl;
  wire[7:0] while_if_mux_12_nl;
  wire[2:0] while_if_mux_13_nl;
  wire[2:0] while_if_mux_14_nl;
  wire while_if_mux_15_nl;

  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_20_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4, rva_in_PopNB_mioi_bcwt);
  assign while_if_mux_1_nl = MUX_v_3_2_2((rva_in_PopNB_mioi_data_data_rsc_z[98:96]),
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_98_96, rva_in_PopNB_mioi_bcwt);
  assign while_if_mux_11_nl = MUX_v_16_2_2((rva_in_PopNB_mioi_data_data_rsc_z[79:64]),
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_79_64, rva_in_PopNB_mioi_bcwt);
  assign while_if_mux_12_nl = MUX_v_8_2_2((rva_in_PopNB_mioi_data_data_rsc_z[55:48]),
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_55_48, rva_in_PopNB_mioi_bcwt);
  assign while_if_mux_13_nl = MUX_v_3_2_2((rva_in_PopNB_mioi_data_data_rsc_z[34:32]),
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_34_32, rva_in_PopNB_mioi_bcwt);
  assign while_if_mux_14_nl = MUX_v_3_2_2((rva_in_PopNB_mioi_data_data_rsc_z[10:8]),
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_10_8, rva_in_PopNB_mioi_bcwt);
  assign while_if_mux_15_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z[0]),
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_0, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = {while_if_mux_1_nl , while_if_mux_11_nl
      , while_if_mux_12_nl , while_if_mux_13_nl , while_if_mux_14_nl , while_if_mux_15_nl};
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_98_96 <= 3'b000;
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_79_64 <= 16'b0000000000000000;
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_55_48 <= 8'b00000000;
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_34_32 <= 3'b000;
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_10_8 <= 3'b000;
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_0 <= 1'b0;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= 20'b00000000000000000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_98_96 <= rva_in_PopNB_mioi_data_data_rsc_z[98:96];
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_79_64 <= rva_in_PopNB_mioi_data_data_rsc_z[79:64];
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_55_48 <= rva_in_PopNB_mioi_data_data_rsc_z[55:48];
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_34_32 <= rva_in_PopNB_mioi_data_data_rsc_z[34:32];
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_10_8 <= rva_in_PopNB_mioi_data_data_rsc_z[10:8];
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt_0 <= rva_in_PopNB_mioi_data_data_rsc_z[0];
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  NMPRun_wen, NMPRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt,
      rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input NMPRun_wen;
  input NMPRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & NMPRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ NMPRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = NMPRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, RVAOutRun_wen, RVAOutRun_wten,
      rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_RVAOutRun,
      rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  input RVAOutRun_wen;
  input RVAOutRun_wten;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [127:0] rva_out_Push_mioi_m_data_rsc_dat_RVAOutRun;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_RVAOutRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_RVAOutRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_RVAOutRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBModule_RVAOutRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl GBModule_RVAOutRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .RVAOutRun_wen(RVAOutRun_wen),
      .RVAOutRun_wten(RVAOutRun_wten),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_RVAOutRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_RVAOutRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_oswt_pff(rva_out_Push_mioi_oswt_pff)
    );
  GBModule_GBModule_RVAOutRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp GBModule_RVAOutRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi (
  clk, rst, nmp_rva_out_vld, nmp_rva_out_rdy, nmp_rva_out_dat, RVAOutRun_wen, RVAOutRun_wten,
      nmp_rva_out_PopNB_mioi_oswt, nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt, nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt,
      RVAOutRun_wten_pff, nmp_rva_out_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input nmp_rva_out_vld;
  output nmp_rva_out_rdy;
  input [127:0] nmp_rva_out_dat;
  input RVAOutRun_wen;
  input RVAOutRun_wten;
  input nmp_rva_out_PopNB_mioi_oswt;
  output [127:0] nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt;
  output nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt;
  input RVAOutRun_wten_pff;
  input nmp_rva_out_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire nmp_rva_out_PopNB_mioi_biwt;
  wire nmp_rva_out_PopNB_mioi_bdwt;
  wire [127:0] nmp_rva_out_PopNB_mioi_data_data_rsc_z;
  wire nmp_rva_out_PopNB_mioi_return_rsc_z;
  wire nmp_rva_out_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB
      nmp_rva_out_PopNB_mioi (
      .this_vld(nmp_rva_out_vld),
      .this_rdy(nmp_rva_out_rdy),
      .this_dat(nmp_rva_out_dat),
      .data_data_rsc_z(nmp_rva_out_PopNB_mioi_data_data_rsc_z),
      .return_rsc_z(nmp_rva_out_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(nmp_rva_out_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi_nmp_rva_out_PopNB_mio_wait_ctrl
      GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi_nmp_rva_out_PopNB_mio_wait_ctrl_inst
      (
      .RVAOutRun_wen(RVAOutRun_wen),
      .RVAOutRun_wten(RVAOutRun_wten),
      .nmp_rva_out_PopNB_mioi_oswt(nmp_rva_out_PopNB_mioi_oswt),
      .nmp_rva_out_PopNB_mioi_biwt(nmp_rva_out_PopNB_mioi_biwt),
      .nmp_rva_out_PopNB_mioi_bdwt(nmp_rva_out_PopNB_mioi_bdwt),
      .nmp_rva_out_PopNB_mioi_biwt_pff(nmp_rva_out_PopNB_mioi_biwt_iff),
      .RVAOutRun_wten_pff(RVAOutRun_wten_pff),
      .nmp_rva_out_PopNB_mioi_oswt_pff(nmp_rva_out_PopNB_mioi_oswt_pff)
    );
  GBModule_GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi_nmp_rva_out_PopNB_mio_wait_dp
      GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi_nmp_rva_out_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt(nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt),
      .nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt(nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt),
      .nmp_rva_out_PopNB_mioi_biwt(nmp_rva_out_PopNB_mioi_biwt),
      .nmp_rva_out_PopNB_mioi_bdwt(nmp_rva_out_PopNB_mioi_bdwt),
      .nmp_rva_out_PopNB_mioi_data_data_rsc_z(nmp_rva_out_PopNB_mioi_data_data_rsc_z),
      .nmp_rva_out_PopNB_mioi_return_rsc_z(nmp_rva_out_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi (
  clk, rst, gbcore_rva_out_vld, gbcore_rva_out_rdy, gbcore_rva_out_dat, RVAOutRun_wen,
      RVAOutRun_wten, gbcore_rva_out_PopNB_mioi_oswt, gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt,
      gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt, RVAOutRun_wten_pff, gbcore_rva_out_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input gbcore_rva_out_vld;
  output gbcore_rva_out_rdy;
  input [127:0] gbcore_rva_out_dat;
  input RVAOutRun_wen;
  input RVAOutRun_wten;
  input gbcore_rva_out_PopNB_mioi_oswt;
  output [127:0] gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt;
  output gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt;
  input RVAOutRun_wten_pff;
  input gbcore_rva_out_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire gbcore_rva_out_PopNB_mioi_biwt;
  wire gbcore_rva_out_PopNB_mioi_bdwt;
  wire [127:0] gbcore_rva_out_PopNB_mioi_data_data_rsc_z;
  wire gbcore_rva_out_PopNB_mioi_return_rsc_z;
  wire gbcore_rva_out_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB
      gbcore_rva_out_PopNB_mioi (
      .this_vld(gbcore_rva_out_vld),
      .this_rdy(gbcore_rva_out_rdy),
      .this_dat(gbcore_rva_out_dat),
      .data_data_rsc_z(gbcore_rva_out_PopNB_mioi_data_data_rsc_z),
      .return_rsc_z(gbcore_rva_out_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(gbcore_rva_out_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi_gbcore_rva_out_PopNB_mio_wait_ctrl
      GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi_gbcore_rva_out_PopNB_mio_wait_ctrl_inst
      (
      .RVAOutRun_wen(RVAOutRun_wen),
      .RVAOutRun_wten(RVAOutRun_wten),
      .gbcore_rva_out_PopNB_mioi_oswt(gbcore_rva_out_PopNB_mioi_oswt),
      .gbcore_rva_out_PopNB_mioi_biwt(gbcore_rva_out_PopNB_mioi_biwt),
      .gbcore_rva_out_PopNB_mioi_bdwt(gbcore_rva_out_PopNB_mioi_bdwt),
      .gbcore_rva_out_PopNB_mioi_biwt_pff(gbcore_rva_out_PopNB_mioi_biwt_iff),
      .RVAOutRun_wten_pff(RVAOutRun_wten_pff),
      .gbcore_rva_out_PopNB_mioi_oswt_pff(gbcore_rva_out_PopNB_mioi_oswt_pff)
    );
  GBModule_GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi_gbcore_rva_out_PopNB_mio_wait_dp
      GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi_gbcore_rva_out_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt(gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt),
      .gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt(gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt),
      .gbcore_rva_out_PopNB_mioi_biwt(gbcore_rva_out_PopNB_mioi_biwt),
      .gbcore_rva_out_PopNB_mioi_bdwt(gbcore_rva_out_PopNB_mioi_bdwt),
      .gbcore_rva_out_PopNB_mioi_data_data_rsc_z(gbcore_rva_out_PopNB_mioi_data_data_rsc_z),
      .gbcore_rva_out_PopNB_mioi_return_rsc_z(gbcore_rva_out_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_nmp_rva_in_Push_mioi
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_nmp_rva_in_Push_mioi (
  clk, rst, nmp_rva_in_vld, nmp_rva_in_rdy, nmp_rva_in_dat, RVAInRun_wen, nmp_rva_in_Push_mioi_oswt,
      nmp_rva_in_Push_mioi_wen_comp, nmp_rva_in_Push_mioi_m_data_rsc_dat_RVAInRun,
      nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun, nmp_rva_in_Push_mioi_m_wstrb_rsc_dat_RVAInRun,
      nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun, nmp_rva_in_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output nmp_rva_in_vld;
  input nmp_rva_in_rdy;
  output [168:0] nmp_rva_in_dat;
  input RVAInRun_wen;
  input nmp_rva_in_Push_mioi_oswt;
  output nmp_rva_in_Push_mioi_wen_comp;
  input [127:0] nmp_rva_in_Push_mioi_m_data_rsc_dat_RVAInRun;
  input [23:0] nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun;
  input [15:0] nmp_rva_in_Push_mioi_m_wstrb_rsc_dat_RVAInRun;
  input nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun;
  input nmp_rva_in_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire nmp_rva_in_Push_mioi_biwt;
  wire nmp_rva_in_Push_mioi_bdwt;
  wire nmp_rva_in_Push_mioi_bcwt;
  wire [23:0] nmp_rva_in_Push_mioi_m_addr_rsc_dat;
  wire nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct;
  wire nmp_rva_in_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [23:0] nl_GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_dp_inst_nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun;
  assign nl_GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_dp_inst_nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun
      = {4'b1100 , (nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun[19:0])};
  GBModule_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_Push
      nmp_rva_in_Push_mioi (
      .this_vld(nmp_rva_in_vld),
      .this_rdy(nmp_rva_in_rdy),
      .this_dat(nmp_rva_in_dat),
      .m_data_rsc_dat(nmp_rva_in_Push_mioi_m_data_rsc_dat_RVAInRun),
      .m_addr_rsc_dat(nmp_rva_in_Push_mioi_m_addr_rsc_dat),
      .m_wstrb_rsc_dat(nmp_rva_in_Push_mioi_m_wstrb_rsc_dat_RVAInRun),
      .m_rw_rsc_dat(nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun),
      .ccs_ccore_start_rsc_dat(nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct),
      .ccs_ccore_done_sync_vld(nmp_rva_in_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_ctrl GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_ctrl_inst
      (
      .RVAInRun_wen(RVAInRun_wen),
      .nmp_rva_in_Push_mioi_oswt(nmp_rva_in_Push_mioi_oswt),
      .nmp_rva_in_Push_mioi_biwt(nmp_rva_in_Push_mioi_biwt),
      .nmp_rva_in_Push_mioi_bdwt(nmp_rva_in_Push_mioi_bdwt),
      .nmp_rva_in_Push_mioi_bcwt(nmp_rva_in_Push_mioi_bcwt),
      .nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct(nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct),
      .nmp_rva_in_Push_mioi_ccs_ccore_done_sync_vld(nmp_rva_in_Push_mioi_ccs_ccore_done_sync_vld),
      .nmp_rva_in_Push_mioi_oswt_pff(nmp_rva_in_Push_mioi_oswt_pff)
    );
  GBModule_GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_dp GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .nmp_rva_in_Push_mioi_oswt(nmp_rva_in_Push_mioi_oswt),
      .nmp_rva_in_Push_mioi_wen_comp(nmp_rva_in_Push_mioi_wen_comp),
      .nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun(nl_GBModule_RVAInRun_nmp_rva_in_Push_mioi_nmp_rva_in_Push_mio_wait_dp_inst_nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun[23:0]),
      .nmp_rva_in_Push_mioi_biwt(nmp_rva_in_Push_mioi_biwt),
      .nmp_rva_in_Push_mioi_bdwt(nmp_rva_in_Push_mioi_bdwt),
      .nmp_rva_in_Push_mioi_bcwt(nmp_rva_in_Push_mioi_bcwt),
      .nmp_rva_in_Push_mioi_m_addr_rsc_dat(nmp_rva_in_Push_mioi_m_addr_rsc_dat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_gbcore_rva_in_Push_mioi
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_gbcore_rva_in_Push_mioi (
  clk, rst, gbcore_rva_in_vld, gbcore_rva_in_rdy, gbcore_rva_in_dat, RVAInRun_wen,
      gbcore_rva_in_Push_mioi_oswt, gbcore_rva_in_Push_mioi_wen_comp, gbcore_rva_in_Push_mioi_m_data_rsc_dat_RVAInRun,
      gbcore_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun, gbcore_rva_in_Push_mioi_m_wstrb_rsc_dat_RVAInRun,
      gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun, gbcore_rva_in_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output gbcore_rva_in_vld;
  input gbcore_rva_in_rdy;
  output [168:0] gbcore_rva_in_dat;
  input RVAInRun_wen;
  input gbcore_rva_in_Push_mioi_oswt;
  output gbcore_rva_in_Push_mioi_wen_comp;
  input [127:0] gbcore_rva_in_Push_mioi_m_data_rsc_dat_RVAInRun;
  input [23:0] gbcore_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun;
  input [15:0] gbcore_rva_in_Push_mioi_m_wstrb_rsc_dat_RVAInRun;
  input gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun;
  input gbcore_rva_in_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire gbcore_rva_in_Push_mioi_biwt;
  wire gbcore_rva_in_Push_mioi_bdwt;
  wire gbcore_rva_in_Push_mioi_bcwt;
  wire gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct;
  wire gbcore_rva_in_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_Push
      gbcore_rva_in_Push_mioi (
      .this_vld(gbcore_rva_in_vld),
      .this_rdy(gbcore_rva_in_rdy),
      .this_dat(gbcore_rva_in_dat),
      .m_data_rsc_dat(gbcore_rva_in_Push_mioi_m_data_rsc_dat_RVAInRun),
      .m_addr_rsc_dat(gbcore_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun),
      .m_wstrb_rsc_dat(gbcore_rva_in_Push_mioi_m_wstrb_rsc_dat_RVAInRun),
      .m_rw_rsc_dat(gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun),
      .ccs_ccore_start_rsc_dat(gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct),
      .ccs_ccore_done_sync_vld(gbcore_rva_in_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBModule_RVAInRun_gbcore_rva_in_Push_mioi_gbcore_rva_in_Push_mio_wait_ctrl
      GBModule_RVAInRun_gbcore_rva_in_Push_mioi_gbcore_rva_in_Push_mio_wait_ctrl_inst
      (
      .RVAInRun_wen(RVAInRun_wen),
      .gbcore_rva_in_Push_mioi_oswt(gbcore_rva_in_Push_mioi_oswt),
      .gbcore_rva_in_Push_mioi_biwt(gbcore_rva_in_Push_mioi_biwt),
      .gbcore_rva_in_Push_mioi_bdwt(gbcore_rva_in_Push_mioi_bdwt),
      .gbcore_rva_in_Push_mioi_bcwt(gbcore_rva_in_Push_mioi_bcwt),
      .gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct(gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun_sct),
      .gbcore_rva_in_Push_mioi_ccs_ccore_done_sync_vld(gbcore_rva_in_Push_mioi_ccs_ccore_done_sync_vld),
      .gbcore_rva_in_Push_mioi_oswt_pff(gbcore_rva_in_Push_mioi_oswt_pff)
    );
  GBModule_GBModule_RVAInRun_gbcore_rva_in_Push_mioi_gbcore_rva_in_Push_mio_wait_dp
      GBModule_RVAInRun_gbcore_rva_in_Push_mioi_gbcore_rva_in_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .gbcore_rva_in_Push_mioi_oswt(gbcore_rva_in_Push_mioi_oswt),
      .gbcore_rva_in_Push_mioi_wen_comp(gbcore_rva_in_Push_mioi_wen_comp),
      .gbcore_rva_in_Push_mioi_biwt(gbcore_rva_in_Push_mioi_biwt),
      .gbcore_rva_in_Push_mioi_bdwt(gbcore_rva_in_Push_mioi_bdwt),
      .gbcore_rva_in_Push_mioi_bcwt(gbcore_rva_in_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, RVAInRun_wen, RVAInRun_wten, rva_in_PopNB_mioi_oswt,
      rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt,
      rva_in_PopNB_mioi_return_rsc_z_mxwt, rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  input RVAInRun_wen;
  input RVAInRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [23:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output [15:0] rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire [15:0] rva_in_PopNB_mioi_data_wstrb_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_wstrb_rsc_z(rva_in_PopNB_mioi_data_wstrb_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBModule_RVAInRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl GBModule_RVAInRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .RVAInRun_wen(RVAInRun_wen),
      .RVAInRun_wten(RVAInRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  GBModule_GBModule_RVAInRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp GBModule_RVAInRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt(rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_wstrb_rsc_z(rva_in_PopNB_mioi_data_wstrb_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi (
  clk, rst, nmp_large_rsp_vld, nmp_large_rsp_rdy, nmp_large_rsp_dat, GBCoreRun_wen,
      nmp_large_rsp_Push_mioi_oswt, nmp_large_rsp_Push_mioi_wen_comp, nmp_large_rsp_Push_mioi_m_read_vector_data_data_rsc_dat_GBCoreRun,
      nmp_large_rsp_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output nmp_large_rsp_vld;
  input nmp_large_rsp_rdy;
  output [127:0] nmp_large_rsp_dat;
  input GBCoreRun_wen;
  input nmp_large_rsp_Push_mioi_oswt;
  output nmp_large_rsp_Push_mioi_wen_comp;
  input [127:0] nmp_large_rsp_Push_mioi_m_read_vector_data_data_rsc_dat_GBCoreRun;
  input nmp_large_rsp_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire nmp_large_rsp_Push_mioi_biwt;
  wire nmp_large_rsp_Push_mioi_bdwt;
  wire nmp_large_rsp_Push_mioi_bcwt;
  wire nmp_large_rsp_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct;
  wire nmp_large_rsp_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_OutBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_Push
      nmp_large_rsp_Push_mioi (
      .this_vld(nmp_large_rsp_vld),
      .this_rdy(nmp_large_rsp_rdy),
      .this_dat(nmp_large_rsp_dat),
      .m_read_vector_data_data_rsc_dat(nmp_large_rsp_Push_mioi_m_read_vector_data_data_rsc_dat_GBCoreRun),
      .ccs_ccore_start_rsc_dat(nmp_large_rsp_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct),
      .ccs_ccore_done_sync_vld(nmp_large_rsp_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_nmp_large_rsp_Push_mio_wait_ctrl
      GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_nmp_large_rsp_Push_mio_wait_ctrl_inst
      (
      .GBCoreRun_wen(GBCoreRun_wen),
      .nmp_large_rsp_Push_mioi_oswt(nmp_large_rsp_Push_mioi_oswt),
      .nmp_large_rsp_Push_mioi_biwt(nmp_large_rsp_Push_mioi_biwt),
      .nmp_large_rsp_Push_mioi_bdwt(nmp_large_rsp_Push_mioi_bdwt),
      .nmp_large_rsp_Push_mioi_bcwt(nmp_large_rsp_Push_mioi_bcwt),
      .nmp_large_rsp_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct(nmp_large_rsp_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct),
      .nmp_large_rsp_Push_mioi_ccs_ccore_done_sync_vld(nmp_large_rsp_Push_mioi_ccs_ccore_done_sync_vld),
      .nmp_large_rsp_Push_mioi_oswt_pff(nmp_large_rsp_Push_mioi_oswt_pff)
    );
  GBModule_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_nmp_large_rsp_Push_mio_wait_dp
      GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_nmp_large_rsp_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .nmp_large_rsp_Push_mioi_oswt(nmp_large_rsp_Push_mioi_oswt),
      .nmp_large_rsp_Push_mioi_wen_comp(nmp_large_rsp_Push_mioi_wen_comp),
      .nmp_large_rsp_Push_mioi_biwt(nmp_large_rsp_Push_mioi_biwt),
      .nmp_large_rsp_Push_mioi_bdwt(nmp_large_rsp_Push_mioi_bdwt),
      .nmp_large_rsp_Push_mioi_bcwt(nmp_large_rsp_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_rva_out_large_Push_mioi
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_rva_out_large_Push_mioi (
  clk, rst, rva_out_large_vld, rva_out_large_rdy, rva_out_large_dat, GBCoreRun_wen,
      rva_out_large_Push_mioi_oswt, rva_out_large_Push_mioi_wen_comp, rva_out_large_Push_mioi_m_data_rsc_dat_GBCoreRun,
      rva_out_large_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_large_vld;
  input rva_out_large_rdy;
  output [127:0] rva_out_large_dat;
  input GBCoreRun_wen;
  input rva_out_large_Push_mioi_oswt;
  output rva_out_large_Push_mioi_wen_comp;
  input [127:0] rva_out_large_Push_mioi_m_data_rsc_dat_GBCoreRun;
  input rva_out_large_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_large_Push_mioi_biwt;
  wire rva_out_large_Push_mioi_bdwt;
  wire rva_out_large_Push_mioi_bcwt;
  wire rva_out_large_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct;
  wire rva_out_large_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_large_Push_mioi (
      .this_vld(rva_out_large_vld),
      .this_rdy(rva_out_large_rdy),
      .this_dat(rva_out_large_dat),
      .m_data_rsc_dat(rva_out_large_Push_mioi_m_data_rsc_dat_GBCoreRun),
      .ccs_ccore_start_rsc_dat(rva_out_large_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_large_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBCore_GBCoreRun_rva_out_large_Push_mioi_rva_out_large_Push_mio_wait_ctrl
      GBCore_GBCoreRun_rva_out_large_Push_mioi_rva_out_large_Push_mio_wait_ctrl_inst
      (
      .GBCoreRun_wen(GBCoreRun_wen),
      .rva_out_large_Push_mioi_oswt(rva_out_large_Push_mioi_oswt),
      .rva_out_large_Push_mioi_biwt(rva_out_large_Push_mioi_biwt),
      .rva_out_large_Push_mioi_bdwt(rva_out_large_Push_mioi_bdwt),
      .rva_out_large_Push_mioi_bcwt(rva_out_large_Push_mioi_bcwt),
      .rva_out_large_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct(rva_out_large_Push_mioi_ccs_ccore_start_rsc_dat_GBCoreRun_sct),
      .rva_out_large_Push_mioi_ccs_ccore_done_sync_vld(rva_out_large_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_large_Push_mioi_oswt_pff(rva_out_large_Push_mioi_oswt_pff)
    );
  GBModule_GBCore_GBCoreRun_rva_out_large_Push_mioi_rva_out_large_Push_mio_wait_dp
      GBCore_GBCoreRun_rva_out_large_Push_mioi_rva_out_large_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_large_Push_mioi_oswt(rva_out_large_Push_mioi_oswt),
      .rva_out_large_Push_mioi_wen_comp(rva_out_large_Push_mioi_wen_comp),
      .rva_out_large_Push_mioi_biwt(rva_out_large_Push_mioi_biwt),
      .rva_out_large_Push_mioi_bdwt(rva_out_large_Push_mioi_bdwt),
      .rva_out_large_Push_mioi_bcwt(rva_out_large_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_nmp_large_req_PopNB_mioi
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_nmp_large_req_PopNB_mioi (
  clk, rst, nmp_large_req_vld, nmp_large_req_rdy, nmp_large_req_dat, GBCoreRun_wen,
      GBCoreRun_wten, nmp_large_req_PopNB_mioi_oswt, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt,
      nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt, nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt,
      nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt, nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt,
      nmp_large_req_PopNB_mioi_return_rsc_z_mxwt, nmp_large_req_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input nmp_large_req_vld;
  output nmp_large_req_rdy;
  input [154:0] nmp_large_req_dat;
  input GBCoreRun_wen;
  input GBCoreRun_wten;
  input nmp_large_req_PopNB_mioi_oswt;
  output nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt;
  output [1:0] nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt;
  output [7:0] nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt;
  output [15:0] nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt;
  output [127:0] nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt;
  output nmp_large_req_PopNB_mioi_return_rsc_z_mxwt;
  input nmp_large_req_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire nmp_large_req_PopNB_mioi_biwt;
  wire nmp_large_req_PopNB_mioi_bdwt;
  wire nmp_large_req_PopNB_mioi_data_is_write_rsc_z;
  wire [1:0] nmp_large_req_PopNB_mioi_data_memory_index_rsc_z;
  wire [7:0] nmp_large_req_PopNB_mioi_data_vector_index_rsc_z;
  wire [15:0] nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z;
  wire [127:0] nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z;
  wire nmp_large_req_PopNB_mioi_return_rsc_z;
  wire nmp_large_req_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB
      nmp_large_req_PopNB_mioi (
      .this_vld(nmp_large_req_vld),
      .this_rdy(nmp_large_req_rdy),
      .this_dat(nmp_large_req_dat),
      .data_is_write_rsc_z(nmp_large_req_PopNB_mioi_data_is_write_rsc_z),
      .data_memory_index_rsc_z(nmp_large_req_PopNB_mioi_data_memory_index_rsc_z),
      .data_vector_index_rsc_z(nmp_large_req_PopNB_mioi_data_vector_index_rsc_z),
      .data_timestep_index_rsc_z(nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z),
      .data_write_data_data_rsc_z(nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z),
      .return_rsc_z(nmp_large_req_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(nmp_large_req_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBCore_GBCoreRun_nmp_large_req_PopNB_mioi_nmp_large_req_PopNB_mio_wait_ctrl
      GBCore_GBCoreRun_nmp_large_req_PopNB_mioi_nmp_large_req_PopNB_mio_wait_ctrl_inst
      (
      .GBCoreRun_wen(GBCoreRun_wen),
      .GBCoreRun_wten(GBCoreRun_wten),
      .nmp_large_req_PopNB_mioi_oswt(nmp_large_req_PopNB_mioi_oswt),
      .nmp_large_req_PopNB_mioi_biwt(nmp_large_req_PopNB_mioi_biwt),
      .nmp_large_req_PopNB_mioi_bdwt(nmp_large_req_PopNB_mioi_bdwt),
      .nmp_large_req_PopNB_mioi_biwt_pff(nmp_large_req_PopNB_mioi_biwt_iff),
      .nmp_large_req_PopNB_mioi_oswt_pff(nmp_large_req_PopNB_mioi_oswt_pff)
    );
  GBModule_GBCore_GBCoreRun_nmp_large_req_PopNB_mioi_nmp_large_req_PopNB_mio_wait_dp
      GBCore_GBCoreRun_nmp_large_req_PopNB_mioi_nmp_large_req_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_return_rsc_z_mxwt(nmp_large_req_PopNB_mioi_return_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_biwt(nmp_large_req_PopNB_mioi_biwt),
      .nmp_large_req_PopNB_mioi_bdwt(nmp_large_req_PopNB_mioi_bdwt),
      .nmp_large_req_PopNB_mioi_data_is_write_rsc_z(nmp_large_req_PopNB_mioi_data_is_write_rsc_z),
      .nmp_large_req_PopNB_mioi_data_memory_index_rsc_z(nmp_large_req_PopNB_mioi_data_memory_index_rsc_z),
      .nmp_large_req_PopNB_mioi_data_vector_index_rsc_z(nmp_large_req_PopNB_mioi_data_vector_index_rsc_z),
      .nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z(nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z),
      .nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z(nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z),
      .nmp_large_req_PopNB_mioi_return_rsc_z(nmp_large_req_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun_rva_in_large_PopNB_mioi
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun_rva_in_large_PopNB_mioi (
  clk, rst, rva_in_large_vld, rva_in_large_rdy, rva_in_large_dat, GBCoreRun_wen,
      GBCoreRun_wten, rva_in_large_PopNB_mioi_oswt, rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt,
      rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt,
      rva_in_large_PopNB_mioi_return_rsc_z_mxwt, rva_in_large_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_large_vld;
  output rva_in_large_rdy;
  input [168:0] rva_in_large_dat;
  input GBCoreRun_wen;
  input GBCoreRun_wten;
  input rva_in_large_PopNB_mioi_oswt;
  output [127:0] rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_large_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_large_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_large_PopNB_mioi_biwt;
  wire rva_in_large_PopNB_mioi_bdwt;
  wire [127:0] rva_in_large_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_large_PopNB_mioi_data_addr_rsc_z;
  wire [15:0] rva_in_large_PopNB_mioi_data_wstrb_rsc_z;
  wire rva_in_large_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_large_PopNB_mioi_return_rsc_z;
  wire [19:0] rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_large_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_large_PopNB_mioi (
      .this_vld(rva_in_large_vld),
      .this_rdy(rva_in_large_rdy),
      .this_dat(rva_in_large_dat),
      .data_data_rsc_z(rva_in_large_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_large_PopNB_mioi_data_addr_rsc_z),
      .data_wstrb_rsc_z(rva_in_large_PopNB_mioi_data_wstrb_rsc_z),
      .data_rw_rsc_z(rva_in_large_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_large_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_large_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_GBCore_GBCoreRun_rva_in_large_PopNB_mioi_rva_in_large_PopNB_mio_wait_ctrl
      GBCore_GBCoreRun_rva_in_large_PopNB_mioi_rva_in_large_PopNB_mio_wait_ctrl_inst
      (
      .GBCoreRun_wen(GBCoreRun_wen),
      .GBCoreRun_wten(GBCoreRun_wten),
      .rva_in_large_PopNB_mioi_oswt(rva_in_large_PopNB_mioi_oswt),
      .rva_in_large_PopNB_mioi_biwt(rva_in_large_PopNB_mioi_biwt),
      .rva_in_large_PopNB_mioi_bdwt(rva_in_large_PopNB_mioi_bdwt),
      .rva_in_large_PopNB_mioi_biwt_pff(rva_in_large_PopNB_mioi_biwt_iff),
      .rva_in_large_PopNB_mioi_oswt_pff(rva_in_large_PopNB_mioi_oswt_pff)
    );
  GBModule_GBCore_GBCoreRun_rva_in_large_PopNB_mioi_rva_in_large_PopNB_mio_wait_dp
      GBCore_GBCoreRun_rva_in_large_PopNB_mioi_rva_in_large_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_large_PopNB_mioi_return_rsc_z_mxwt(rva_in_large_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_large_PopNB_mioi_biwt(rva_in_large_PopNB_mioi_biwt),
      .rva_in_large_PopNB_mioi_bdwt(rva_in_large_PopNB_mioi_bdwt),
      .rva_in_large_PopNB_mioi_data_data_rsc_z(rva_in_large_PopNB_mioi_data_data_rsc_z),
      .rva_in_large_PopNB_mioi_data_addr_rsc_z(rva_in_large_PopNB_mioi_data_addr_rsc_z),
      .rva_in_large_PopNB_mioi_data_rw_rsc_z(rva_in_large_PopNB_mioi_data_rw_rsc_z),
      .rva_in_large_PopNB_mioi_return_rsc_z(rva_in_large_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_done_Push_mioi
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_done_Push_mioi (
  clk, rst, done_vld, done_rdy, done_dat, NMPRun_wen, done_Push_mioi_oswt, done_Push_mioi_wen_comp,
      done_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output done_vld;
  input done_rdy;
  output done_dat;
  input NMPRun_wen;
  input done_Push_mioi_oswt;
  output done_Push_mioi_wen_comp;
  input done_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire done_Push_mioi_biwt;
  wire done_Push_mioi_bdwt;
  wire done_Push_mioi_bcwt;
  wire done_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct;
  wire done_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_OutBlocking_bool_Connections_SYN_PORT_Push  done_Push_mioi
      (
      .this_vld(done_vld),
      .this_rdy(done_rdy),
      .this_dat(done_dat),
      .ccs_ccore_start_rsc_dat(done_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct),
      .ccs_ccore_done_sync_vld(done_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_NMP_NMPRun_done_Push_mioi_done_Push_mio_wait_ctrl NMP_NMPRun_done_Push_mioi_done_Push_mio_wait_ctrl_inst
      (
      .NMPRun_wen(NMPRun_wen),
      .done_Push_mioi_oswt(done_Push_mioi_oswt),
      .done_Push_mioi_biwt(done_Push_mioi_biwt),
      .done_Push_mioi_bdwt(done_Push_mioi_bdwt),
      .done_Push_mioi_bcwt(done_Push_mioi_bcwt),
      .done_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct(done_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct),
      .done_Push_mioi_ccs_ccore_done_sync_vld(done_Push_mioi_ccs_ccore_done_sync_vld),
      .done_Push_mioi_oswt_pff(done_Push_mioi_oswt_pff)
    );
  GBModule_NMP_NMPRun_done_Push_mioi_done_Push_mio_wait_dp NMP_NMPRun_done_Push_mioi_done_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_Push_mioi_oswt(done_Push_mioi_oswt),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp),
      .done_Push_mioi_biwt(done_Push_mioi_biwt),
      .done_Push_mioi_bdwt(done_Push_mioi_bdwt),
      .done_Push_mioi_bcwt(done_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, NMPRun_wen, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff, rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  input NMPRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [127:0] rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire [127:0] rva_out_Push_mioi_m_data_rsc_dat;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [127:0] nl_NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst_rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff;
  assign nl_NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst_rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff
      = {29'b00000000000000000000000000000 , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[98:96])
      , 16'b0000000000000000 , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[79:64])
      , 8'b00000000 , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[55:48]) , 13'b0000000000000
      , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[34:32]) , 21'b000000000000000000000
      , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[10:8]) , 7'b0000000 , (rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[0])};
  GBModule_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .NMPRun_wen(NMPRun_wen),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_NMPRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_oswt_pff(rva_out_Push_mioi_oswt_pff)
    );
  GBModule_NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat),
      .rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff(nl_NMP_NMPRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst_rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[127:0])
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_large_rsp_PopNB_mioi
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_large_rsp_PopNB_mioi (
  clk, rst, large_rsp_vld, large_rsp_rdy, large_rsp_dat, NMPRun_wen, NMPRun_wten,
      large_rsp_PopNB_mioi_oswt, large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt,
      large_rsp_PopNB_mioi_return_rsc_z_mxwt, large_rsp_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input large_rsp_vld;
  output large_rsp_rdy;
  input [127:0] large_rsp_dat;
  input NMPRun_wen;
  input NMPRun_wten;
  input large_rsp_PopNB_mioi_oswt;
  output [127:0] large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt;
  output large_rsp_PopNB_mioi_return_rsc_z_mxwt;
  input large_rsp_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire large_rsp_PopNB_mioi_biwt;
  wire large_rsp_PopNB_mioi_bdwt;
  wire [127:0] large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z;
  wire large_rsp_PopNB_mioi_return_rsc_z;
  wire large_rsp_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_InBlocking_spec_GB_Large_DataRsp_1U_Connections_SYN_PORT_PopNB
      large_rsp_PopNB_mioi (
      .this_vld(large_rsp_vld),
      .this_rdy(large_rsp_rdy),
      .this_dat(large_rsp_dat),
      .data_read_vector_data_data_rsc_z(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z),
      .return_rsc_z(large_rsp_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(large_rsp_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_NMP_NMPRun_large_rsp_PopNB_mioi_large_rsp_PopNB_mio_wait_ctrl NMP_NMPRun_large_rsp_PopNB_mioi_large_rsp_PopNB_mio_wait_ctrl_inst
      (
      .NMPRun_wen(NMPRun_wen),
      .NMPRun_wten(NMPRun_wten),
      .large_rsp_PopNB_mioi_oswt(large_rsp_PopNB_mioi_oswt),
      .large_rsp_PopNB_mioi_biwt(large_rsp_PopNB_mioi_biwt),
      .large_rsp_PopNB_mioi_bdwt(large_rsp_PopNB_mioi_bdwt),
      .large_rsp_PopNB_mioi_biwt_pff(large_rsp_PopNB_mioi_biwt_iff),
      .large_rsp_PopNB_mioi_oswt_pff(large_rsp_PopNB_mioi_oswt_pff)
    );
  GBModule_NMP_NMPRun_large_rsp_PopNB_mioi_large_rsp_PopNB_mio_wait_dp NMP_NMPRun_large_rsp_PopNB_mioi_large_rsp_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt),
      .large_rsp_PopNB_mioi_return_rsc_z_mxwt(large_rsp_PopNB_mioi_return_rsc_z_mxwt),
      .large_rsp_PopNB_mioi_biwt(large_rsp_PopNB_mioi_biwt),
      .large_rsp_PopNB_mioi_bdwt(large_rsp_PopNB_mioi_bdwt),
      .large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z),
      .large_rsp_PopNB_mioi_return_rsc_z(large_rsp_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_start_PopNB_mioi
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_start_PopNB_mioi (
  clk, rst, start_vld, start_rdy, start_dat, NMPRun_wen, NMPRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input NMPRun_wen;
  input NMPRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_vld(start_vld),
      .this_rdy(start_rdy),
      .this_dat(start_dat),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_NMP_NMPRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl NMP_NMPRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .NMPRun_wen(NMPRun_wen),
      .NMPRun_wten(NMPRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_biwt_pff(start_PopNB_mioi_biwt_iff),
      .start_PopNB_mioi_oswt_pff(start_PopNB_mioi_oswt_pff)
    );
  GBModule_NMP_NMPRun_start_PopNB_mioi_start_PopNB_mio_wait_dp NMP_NMPRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_large_req_Push_mioi
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_large_req_Push_mioi (
  clk, rst, large_req_vld, large_req_rdy, large_req_dat, NMPRun_wen, large_req_Push_mioi_oswt,
      large_req_Push_mioi_wen_comp, large_req_Push_mioi_m_is_write_rsc_dat_NMPRun,
      large_req_Push_mioi_m_memory_index_rsc_dat_NMPRun, large_req_Push_mioi_m_vector_index_rsc_dat_NMPRun,
      large_req_Push_mioi_m_timestep_index_rsc_dat_NMPRun, large_req_Push_mioi_m_write_data_data_rsc_dat_NMPRun,
      large_req_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output large_req_vld;
  input large_req_rdy;
  output [154:0] large_req_dat;
  input NMPRun_wen;
  input large_req_Push_mioi_oswt;
  output large_req_Push_mioi_wen_comp;
  input large_req_Push_mioi_m_is_write_rsc_dat_NMPRun;
  input [1:0] large_req_Push_mioi_m_memory_index_rsc_dat_NMPRun;
  input [7:0] large_req_Push_mioi_m_vector_index_rsc_dat_NMPRun;
  input [15:0] large_req_Push_mioi_m_timestep_index_rsc_dat_NMPRun;
  input [127:0] large_req_Push_mioi_m_write_data_data_rsc_dat_NMPRun;
  input large_req_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire large_req_Push_mioi_biwt;
  wire large_req_Push_mioi_bdwt;
  wire large_req_Push_mioi_bcwt;
  wire large_req_Push_mioi_m_is_write_rsc_dat_NMPRun_sct;
  wire large_req_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_OutBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_Push
      large_req_Push_mioi (
      .this_vld(large_req_vld),
      .this_rdy(large_req_rdy),
      .this_dat(large_req_dat),
      .m_is_write_rsc_dat(large_req_Push_mioi_m_is_write_rsc_dat_NMPRun),
      .m_memory_index_rsc_dat(large_req_Push_mioi_m_memory_index_rsc_dat_NMPRun),
      .m_vector_index_rsc_dat(large_req_Push_mioi_m_vector_index_rsc_dat_NMPRun),
      .m_timestep_index_rsc_dat(large_req_Push_mioi_m_timestep_index_rsc_dat_NMPRun),
      .m_write_data_data_rsc_dat(large_req_Push_mioi_m_write_data_data_rsc_dat_NMPRun),
      .ccs_ccore_start_rsc_dat(large_req_Push_mioi_m_is_write_rsc_dat_NMPRun_sct),
      .ccs_ccore_done_sync_vld(large_req_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_NMP_NMPRun_large_req_Push_mioi_large_req_Push_mio_wait_ctrl NMP_NMPRun_large_req_Push_mioi_large_req_Push_mio_wait_ctrl_inst
      (
      .NMPRun_wen(NMPRun_wen),
      .large_req_Push_mioi_oswt(large_req_Push_mioi_oswt),
      .large_req_Push_mioi_biwt(large_req_Push_mioi_biwt),
      .large_req_Push_mioi_bdwt(large_req_Push_mioi_bdwt),
      .large_req_Push_mioi_bcwt(large_req_Push_mioi_bcwt),
      .large_req_Push_mioi_m_is_write_rsc_dat_NMPRun_sct(large_req_Push_mioi_m_is_write_rsc_dat_NMPRun_sct),
      .large_req_Push_mioi_ccs_ccore_done_sync_vld(large_req_Push_mioi_ccs_ccore_done_sync_vld),
      .large_req_Push_mioi_oswt_pff(large_req_Push_mioi_oswt_pff)
    );
  GBModule_NMP_NMPRun_large_req_Push_mioi_large_req_Push_mio_wait_dp NMP_NMPRun_large_req_Push_mioi_large_req_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .large_req_Push_mioi_oswt(large_req_Push_mioi_oswt),
      .large_req_Push_mioi_wen_comp(large_req_Push_mioi_wen_comp),
      .large_req_Push_mioi_biwt(large_req_Push_mioi_biwt),
      .large_req_Push_mioi_bdwt(large_req_Push_mioi_bdwt),
      .large_req_Push_mioi_bcwt(large_req_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, NMPRun_wen, NMPRun_wten, rva_in_PopNB_mioi_oswt,
      rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  input NMPRun_wen;
  input NMPRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [33:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire [15:0] rva_in_PopNB_mioi_data_wstrb_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire [33:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt_pconst;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_wstrb_rsc_z(rva_in_PopNB_mioi_data_wstrb_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  GBModule_NMP_NMPRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl NMP_NMPRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .NMPRun_wen(NMPRun_wen),
      .NMPRun_wten(NMPRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  GBModule_NMP_NMPRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp NMP_NMPRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = rva_in_PopNB_mioi_data_data_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAOutRun
// ------------------------------------------------------------------


module GBModule_GBModule_RVAOutRun (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, gbcore_rva_out_vld, gbcore_rva_out_rdy,
      gbcore_rva_out_dat, nmp_rva_out_vld, nmp_rva_out_rdy, nmp_rva_out_dat
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  input gbcore_rva_out_vld;
  output gbcore_rva_out_rdy;
  input [127:0] gbcore_rva_out_dat;
  input nmp_rva_out_vld;
  output nmp_rva_out_rdy;
  input [127:0] nmp_rva_out_dat;


  // Interconnect Declarations
  wire RVAOutRun_wten;
  wire [127:0] gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt;
  wire gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt;
  wire [127:0] nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt;
  wire nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire fsm_output;
  reg while_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB_return_sva_1;
  reg while_stage_0_3;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_nmp_rva_out_PopNB_mioi_iswt0_cse;
  reg reg_gbcore_rva_out_PopNB_mioi_iswt0_cse;
  wire RVAOutRun_wten_iff;
  wire and_3_rmff;
  wire and_2_rmff;
  reg [127:0] while_rva_out_reg_data_sva_1;


  // Interconnect Declarations for Component Instantiations 
  wire and_1_nl;
  wire [127:0] nl_GBModule_RVAOutRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_RVAOutRun;
  assign and_1_nl = fsm_output & (~ while_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nl_GBModule_RVAOutRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_RVAOutRun
      = MUX_v_128_2_2(while_rva_out_reg_data_sva_1, nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt,
      and_1_nl);
  GBModule_GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi GBModule_RVAOutRun_gbcore_rva_out_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .gbcore_rva_out_vld(gbcore_rva_out_vld),
      .gbcore_rva_out_rdy(gbcore_rva_out_rdy),
      .gbcore_rva_out_dat(gbcore_rva_out_dat),
      .RVAOutRun_wen(rva_out_Push_mioi_wen_comp),
      .RVAOutRun_wten(RVAOutRun_wten),
      .gbcore_rva_out_PopNB_mioi_oswt(reg_gbcore_rva_out_PopNB_mioi_iswt0_cse),
      .gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt(gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt),
      .gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt(gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt),
      .RVAOutRun_wten_pff(RVAOutRun_wten_iff),
      .gbcore_rva_out_PopNB_mioi_oswt_pff(fsm_output)
    );
  GBModule_GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi GBModule_RVAOutRun_nmp_rva_out_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .nmp_rva_out_vld(nmp_rva_out_vld),
      .nmp_rva_out_rdy(nmp_rva_out_rdy),
      .nmp_rva_out_dat(nmp_rva_out_dat),
      .RVAOutRun_wen(rva_out_Push_mioi_wen_comp),
      .RVAOutRun_wten(RVAOutRun_wten),
      .nmp_rva_out_PopNB_mioi_oswt(reg_nmp_rva_out_PopNB_mioi_iswt0_cse),
      .nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt(nmp_rva_out_PopNB_mioi_data_data_rsc_z_mxwt),
      .nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt(nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt),
      .RVAOutRun_wten_pff(RVAOutRun_wten_iff),
      .nmp_rva_out_PopNB_mioi_oswt_pff(and_3_rmff)
    );
  GBModule_GBModule_RVAOutRun_rva_out_Push_mioi GBModule_RVAOutRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .RVAOutRun_wen(rva_out_Push_mioi_wen_comp),
      .RVAOutRun_wten(RVAOutRun_wten_iff),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_RVAOutRun(nl_GBModule_RVAOutRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_RVAOutRun[127:0]),
      .rva_out_Push_mioi_oswt_pff(and_2_rmff)
    );
  GBModule_GBModule_RVAOutRun_staller_1 GBModule_RVAOutRun_staller_1_inst (
      .clk(clk),
      .rst(rst),
      .RVAOutRun_wten(RVAOutRun_wten),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .RVAOutRun_wten_pff(RVAOutRun_wten_iff)
    );
  GBModule_GBModule_RVAOutRun_RVAOutRun_fsm GBModule_RVAOutRun_RVAOutRun_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .fsm_output(fsm_output)
    );
  assign and_2_rmff = (nmp_rva_out_PopNB_mioi_return_rsc_z_mxwt | while_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign and_3_rmff = reg_gbcore_rva_out_PopNB_mioi_iswt0_cse & (~ gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_nmp_rva_out_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_gbcore_rva_out_PopNB_mioi_iswt0_cse <= 1'b0;
      while_stage_0_3 <= 1'b0;
    end
    else if ( rva_out_Push_mioi_wen_comp ) begin
      reg_rva_out_Push_mioi_iswt0_cse <= and_2_rmff;
      reg_nmp_rva_out_PopNB_mioi_iswt0_cse <= and_3_rmff;
      reg_gbcore_rva_out_PopNB_mioi_iswt0_cse <= fsm_output;
      while_stage_0_3 <= reg_gbcore_rva_out_PopNB_mioi_iswt0_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB_return_sva_1
          <= 1'b0;
    end
    else if ( rva_out_Push_mioi_wen_comp & reg_gbcore_rva_out_PopNB_mioi_iswt0_cse
        ) begin
      while_Connections_Combinational_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_PopNB_return_sva_1
          <= gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_rva_out_reg_data_sva_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rva_out_Push_mioi_wen_comp & reg_gbcore_rva_out_PopNB_mioi_iswt0_cse
        & gbcore_rva_out_PopNB_mioi_return_rsc_z_mxwt ) begin
      while_rva_out_reg_data_sva_1 <= gbcore_rva_out_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBModule_RVAInRun
// ------------------------------------------------------------------


module GBModule_GBModule_RVAInRun (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, gbcore_rva_in_vld, gbcore_rva_in_rdy,
      gbcore_rva_in_dat, nmp_rva_in_vld, nmp_rva_in_rdy, nmp_rva_in_dat, SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output gbcore_rva_in_vld;
  input gbcore_rva_in_rdy;
  output [168:0] gbcore_rva_in_dat;
  output nmp_rva_in_vld;
  input nmp_rva_in_rdy;
  output [168:0] nmp_rva_in_dat;
  output [31:0] SC_SRAM_CONFIG;
  reg [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire RVAInRun_wen;
  wire RVAInRun_wten;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire [15:0] rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire gbcore_rva_in_Push_mioi_wen_comp;
  wire nmp_rva_in_Push_mioi_wen_comp;
  wire fsm_output;
  wire and_dcpl_2;
  reg reg_nmp_rva_in_Push_mioi_iswt0_cse;
  reg reg_gbcore_rva_in_Push_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire and_6_rmff;
  wire and_4_rmff;

  wire mux_1_nl;
  wire mux_nl;
  wire nor_nl;
  wire or_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [23:0] nl_GBModule_RVAInRun_nmp_rva_in_Push_mioi_inst_nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun;
  assign nl_GBModule_RVAInRun_nmp_rva_in_Push_mioi_inst_nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun
      = {4'b1100 , (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:0])};
  GBModule_GBModule_RVAInRun_rva_in_PopNB_mioi GBModule_RVAInRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .RVAInRun_wen(RVAInRun_wen),
      .RVAInRun_wten(RVAInRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt(rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(fsm_output)
    );
  GBModule_GBModule_RVAInRun_gbcore_rva_in_Push_mioi GBModule_RVAInRun_gbcore_rva_in_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .gbcore_rva_in_vld(gbcore_rva_in_vld),
      .gbcore_rva_in_rdy(gbcore_rva_in_rdy),
      .gbcore_rva_in_dat(gbcore_rva_in_dat),
      .RVAInRun_wen(RVAInRun_wen),
      .gbcore_rva_in_Push_mioi_oswt(reg_gbcore_rva_in_Push_mioi_iswt0_cse),
      .gbcore_rva_in_Push_mioi_wen_comp(gbcore_rva_in_Push_mioi_wen_comp),
      .gbcore_rva_in_Push_mioi_m_data_rsc_dat_RVAInRun(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .gbcore_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .gbcore_rva_in_Push_mioi_m_wstrb_rsc_dat_RVAInRun(rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt),
      .gbcore_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .gbcore_rva_in_Push_mioi_oswt_pff(and_6_rmff)
    );
  GBModule_GBModule_RVAInRun_nmp_rva_in_Push_mioi GBModule_RVAInRun_nmp_rva_in_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .nmp_rva_in_vld(nmp_rva_in_vld),
      .nmp_rva_in_rdy(nmp_rva_in_rdy),
      .nmp_rva_in_dat(nmp_rva_in_dat),
      .RVAInRun_wen(RVAInRun_wen),
      .nmp_rva_in_Push_mioi_oswt(reg_nmp_rva_in_Push_mioi_iswt0_cse),
      .nmp_rva_in_Push_mioi_wen_comp(nmp_rva_in_Push_mioi_wen_comp),
      .nmp_rva_in_Push_mioi_m_data_rsc_dat_RVAInRun(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun(nl_GBModule_RVAInRun_nmp_rva_in_Push_mioi_inst_nmp_rva_in_Push_mioi_m_addr_rsc_dat_RVAInRun[23:0]),
      .nmp_rva_in_Push_mioi_m_wstrb_rsc_dat_RVAInRun(rva_in_PopNB_mioi_data_wstrb_rsc_z_mxwt),
      .nmp_rva_in_Push_mioi_m_rw_rsc_dat_RVAInRun(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .nmp_rva_in_Push_mioi_oswt_pff(and_4_rmff)
    );
  GBModule_GBModule_RVAInRun_staller GBModule_RVAInRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .RVAInRun_wen(RVAInRun_wen),
      .RVAInRun_wten(RVAInRun_wten),
      .gbcore_rva_in_Push_mioi_wen_comp(gbcore_rva_in_Push_mioi_wen_comp),
      .nmp_rva_in_Push_mioi_wen_comp(nmp_rva_in_Push_mioi_wen_comp)
    );
  GBModule_GBModule_RVAInRun_RVAInRun_fsm GBModule_RVAInRun_RVAInRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .RVAInRun_wen(RVAInRun_wen),
      .fsm_output(fsm_output)
    );
  assign and_4_rmff = and_dcpl_2 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[23:20]==4'b1100);
  assign mux_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[21]), (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[21])),
      rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[22]);
  assign nor_nl = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[22:21]!=2'b10));
  assign or_nl = (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[20])) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign mux_1_nl = MUX_s_1_2_2(mux_nl, nor_nl, or_nl);
  assign and_6_rmff = mux_1_nl & and_dcpl_2 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[23]));
  assign and_dcpl_2 = reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nmp_rva_in_Push_mioi_iswt0_cse <= 1'b0;
      reg_gbcore_rva_in_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
    end
    else if ( RVAInRun_wen ) begin
      reg_nmp_rva_in_Push_mioi_iswt0_cse <= and_4_rmff;
      reg_gbcore_rva_in_Push_mioi_iswt0_cse <= and_6_rmff;
      reg_rva_in_PopNB_mioi_iswt0_cse <= fsm_output;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      SC_SRAM_CONFIG <= 32'b00000000000000000000000000000000;
    end
    else if ( RVAInRun_wen & (~((~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_return_rsc_z_mxwt))
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[22:21]!=2'b01) | (~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[20]))) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[23])))
        ) begin
      SC_SRAM_CONFIG <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:0];
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore_GBCoreRun
// ------------------------------------------------------------------


module GBModule_GBCore_GBCoreRun (
  clk, rst, rva_in_large_vld, rva_in_large_rdy, rva_in_large_dat, rva_out_large_vld,
      rva_out_large_rdy, rva_out_large_dat, nmp_large_req_vld, nmp_large_req_rdy,
      nmp_large_req_dat, nmp_large_rsp_vld, nmp_large_rsp_rdy, nmp_large_rsp_dat,
      SC_SRAM_CONFIG, large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d, large_mem_banks_bank_a0_a0_a0_a0_a_rsci_d_d,
      large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d, large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d,
      large_mem_banks_bank_a0_a0_a0_a1_a_rsci_d_d, large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d,
      large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d, large_mem_banks_bank_a0_a0_a1_a0_a_rsci_d_d,
      large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d, large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d,
      large_mem_banks_bank_a0_a0_a1_a1_a_rsci_d_d, large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d,
      large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d, large_mem_banks_bank_a0_a1_a0_a0_a_rsci_d_d,
      large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d, large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d,
      large_mem_banks_bank_a0_a1_a0_a1_a_rsci_d_d, large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d,
      large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d, large_mem_banks_bank_a0_a1_a1_a0_a_rsci_d_d,
      large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d, large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d,
      large_mem_banks_bank_a0_a1_a1_a1_a_rsci_d_d, large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d,
      large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d, large_mem_banks_bank_a1_a0_a0_a0_a_rsci_d_d,
      large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d, large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d,
      large_mem_banks_bank_a1_a0_a0_a1_a_rsci_d_d, large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d,
      large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d, large_mem_banks_bank_a1_a0_a1_a0_a_rsci_d_d,
      large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d, large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d,
      large_mem_banks_bank_a1_a0_a1_a1_a_rsci_d_d, large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d,
      large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d, large_mem_banks_bank_a1_a1_a0_a0_a_rsci_d_d,
      large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d, large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d,
      large_mem_banks_bank_a1_a1_a0_a1_a_rsci_d_d, large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d,
      large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d, large_mem_banks_bank_a1_a1_a1_a0_a_rsci_d_d,
      large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d, large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d,
      large_mem_banks_bank_a1_a1_a1_a1_a_rsci_d_d, large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d,
      GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_a, GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_b,
      GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_c, GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_z,
      large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_pff, large_mem_banks_bank_a0_a0_a0_a0_a_rsci_re_d_pff,
      large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_pff, large_mem_banks_bank_a0_a0_a0_a0_a_rsci_we_d_pff,
      large_mem_banks_bank_a0_a0_a0_a1_a_rsci_re_d_pff, large_mem_banks_bank_a0_a0_a0_a1_a_rsci_we_d_pff,
      large_mem_banks_bank_a0_a0_a1_a0_a_rsci_re_d_pff, large_mem_banks_bank_a0_a0_a1_a0_a_rsci_we_d_pff,
      large_mem_banks_bank_a0_a0_a1_a1_a_rsci_re_d_pff, large_mem_banks_bank_a0_a0_a1_a1_a_rsci_we_d_pff,
      large_mem_banks_bank_a0_a1_a0_a0_a_rsci_re_d_pff, large_mem_banks_bank_a0_a1_a0_a0_a_rsci_we_d_pff,
      large_mem_banks_bank_a0_a1_a0_a1_a_rsci_re_d_pff, large_mem_banks_bank_a0_a1_a0_a1_a_rsci_we_d_pff,
      large_mem_banks_bank_a0_a1_a1_a0_a_rsci_re_d_pff, large_mem_banks_bank_a0_a1_a1_a0_a_rsci_we_d_pff,
      large_mem_banks_bank_a0_a1_a1_a1_a_rsci_re_d_pff, large_mem_banks_bank_a0_a1_a1_a1_a_rsci_we_d_pff,
      large_mem_banks_bank_a1_a0_a0_a0_a_rsci_re_d_pff, large_mem_banks_bank_a1_a0_a0_a0_a_rsci_we_d_pff,
      large_mem_banks_bank_a1_a0_a0_a1_a_rsci_re_d_pff, large_mem_banks_bank_a1_a0_a0_a1_a_rsci_we_d_pff,
      large_mem_banks_bank_a1_a0_a1_a0_a_rsci_re_d_pff, large_mem_banks_bank_a1_a0_a1_a0_a_rsci_we_d_pff,
      large_mem_banks_bank_a1_a0_a1_a1_a_rsci_re_d_pff, large_mem_banks_bank_a1_a0_a1_a1_a_rsci_we_d_pff,
      large_mem_banks_bank_a1_a1_a0_a0_a_rsci_re_d_pff, large_mem_banks_bank_a1_a1_a0_a0_a_rsci_we_d_pff,
      large_mem_banks_bank_a1_a1_a0_a1_a_rsci_re_d_pff, large_mem_banks_bank_a1_a1_a0_a1_a_rsci_we_d_pff,
      large_mem_banks_bank_a1_a1_a1_a0_a_rsci_re_d_pff, large_mem_banks_bank_a1_a1_a1_a0_a_rsci_we_d_pff,
      large_mem_banks_bank_a1_a1_a1_a1_a_rsci_re_d_pff, large_mem_banks_bank_a1_a1_a1_a1_a_rsci_we_d_pff
);
  input clk;
  input rst;
  input rva_in_large_vld;
  output rva_in_large_rdy;
  input [168:0] rva_in_large_dat;
  output rva_out_large_vld;
  input rva_out_large_rdy;
  output [127:0] rva_out_large_dat;
  input nmp_large_req_vld;
  output nmp_large_req_rdy;
  input [154:0] nmp_large_req_dat;
  output nmp_large_rsp_vld;
  input nmp_large_rsp_rdy;
  output [127:0] nmp_large_rsp_dat;
  input [31:0] SC_SRAM_CONFIG;
  output large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d;
  output large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a0_a0_a0_a1_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d;
  output large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a0_a0_a1_a0_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d;
  output large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a0_a0_a1_a1_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d;
  output large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a0_a1_a0_a0_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d;
  output large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a0_a1_a0_a1_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d;
  output large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a0_a1_a1_a0_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d;
  output large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a0_a1_a1_a1_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d;
  output large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a1_a0_a0_a0_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d;
  output large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a1_a0_a0_a1_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d;
  output large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a1_a0_a1_a0_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d;
  output large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a1_a0_a1_a1_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d;
  output large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a1_a1_a0_a0_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d;
  output large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a1_a1_a0_a1_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d;
  output large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a1_a1_a1_a0_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d;
  output large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d;
  output [127:0] large_mem_banks_bank_a1_a1_a1_a1_a_rsci_d_d;
  input [127:0] large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d;
  output [7:0] GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_a;
  output [15:0] GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_b;
  output [11:0] GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_c;
  input [15:0] GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_z;
  output [11:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_pff;
  output large_mem_banks_bank_a0_a0_a0_a0_a_rsci_re_d_pff;
  output [11:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_pff;
  output large_mem_banks_bank_a0_a0_a0_a0_a_rsci_we_d_pff;
  output large_mem_banks_bank_a0_a0_a0_a1_a_rsci_re_d_pff;
  output large_mem_banks_bank_a0_a0_a0_a1_a_rsci_we_d_pff;
  output large_mem_banks_bank_a0_a0_a1_a0_a_rsci_re_d_pff;
  output large_mem_banks_bank_a0_a0_a1_a0_a_rsci_we_d_pff;
  output large_mem_banks_bank_a0_a0_a1_a1_a_rsci_re_d_pff;
  output large_mem_banks_bank_a0_a0_a1_a1_a_rsci_we_d_pff;
  output large_mem_banks_bank_a0_a1_a0_a0_a_rsci_re_d_pff;
  output large_mem_banks_bank_a0_a1_a0_a0_a_rsci_we_d_pff;
  output large_mem_banks_bank_a0_a1_a0_a1_a_rsci_re_d_pff;
  output large_mem_banks_bank_a0_a1_a0_a1_a_rsci_we_d_pff;
  output large_mem_banks_bank_a0_a1_a1_a0_a_rsci_re_d_pff;
  output large_mem_banks_bank_a0_a1_a1_a0_a_rsci_we_d_pff;
  output large_mem_banks_bank_a0_a1_a1_a1_a_rsci_re_d_pff;
  output large_mem_banks_bank_a0_a1_a1_a1_a_rsci_we_d_pff;
  output large_mem_banks_bank_a1_a0_a0_a0_a_rsci_re_d_pff;
  output large_mem_banks_bank_a1_a0_a0_a0_a_rsci_we_d_pff;
  output large_mem_banks_bank_a1_a0_a0_a1_a_rsci_re_d_pff;
  output large_mem_banks_bank_a1_a0_a0_a1_a_rsci_we_d_pff;
  output large_mem_banks_bank_a1_a0_a1_a0_a_rsci_re_d_pff;
  output large_mem_banks_bank_a1_a0_a1_a0_a_rsci_we_d_pff;
  output large_mem_banks_bank_a1_a0_a1_a1_a_rsci_re_d_pff;
  output large_mem_banks_bank_a1_a0_a1_a1_a_rsci_we_d_pff;
  output large_mem_banks_bank_a1_a1_a0_a0_a_rsci_re_d_pff;
  output large_mem_banks_bank_a1_a1_a0_a0_a_rsci_we_d_pff;
  output large_mem_banks_bank_a1_a1_a0_a1_a_rsci_re_d_pff;
  output large_mem_banks_bank_a1_a1_a0_a1_a_rsci_we_d_pff;
  output large_mem_banks_bank_a1_a1_a1_a0_a_rsci_re_d_pff;
  output large_mem_banks_bank_a1_a1_a1_a0_a_rsci_we_d_pff;
  output large_mem_banks_bank_a1_a1_a1_a1_a_rsci_re_d_pff;
  output large_mem_banks_bank_a1_a1_a1_a1_a_rsci_we_d_pff;


  // Interconnect Declarations
  wire GBCoreRun_wen;
  wire GBCoreRun_wten;
  wire [127:0] rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [19:0] rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_large_PopNB_mioi_return_rsc_z_mxwt;
  wire nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt;
  wire [1:0] nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt;
  wire [7:0] nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt;
  wire [15:0] nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt;
  wire [127:0] nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt;
  wire nmp_large_req_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_large_Push_mioi_wen_comp;
  wire nmp_large_rsp_Push_mioi_wen_comp;
  wire fsm_output;
  wire [15:0] large_mem_write_arbxbar_xbar_for_lshift_tmp;
  wire [15:0] large_mem_read_arbxbar_xbar_for_1_lshift_tmp;
  wire crossbar_spec_GB_Large_WordType_16U_16U_for_mux_tmp;
  wire large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_and_tmp;
  wire [2:0] while_mux_2_tmp;
  wire and_dcpl_1;
  wire or_dcpl_1;
  wire and_dcpl_7;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_10;
  wire and_dcpl_11;
  wire and_dcpl_12;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire and_dcpl_17;
  wire and_dcpl_18;
  wire and_dcpl_19;
  wire and_dcpl_20;
  wire and_dcpl_21;
  wire and_dcpl_22;
  wire and_dcpl_24;
  wire and_dcpl_26;
  wire and_dcpl_28;
  wire and_dcpl_30;
  wire and_dcpl_32;
  wire and_dcpl_34;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire and_dcpl_40;
  wire and_dcpl_42;
  wire and_dcpl_44;
  wire and_dcpl_46;
  wire and_dcpl_48;
  wire and_dcpl_50;
  wire and_dcpl_52;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_63;
  wire and_dcpl_72;
  wire or_tmp_11;
  wire and_dcpl_93;
  wire and_dcpl_94;
  wire and_dcpl_95;
  wire and_dcpl_199;
  wire and_dcpl_204;
  wire and_dcpl_206;
  wire or_dcpl_71;
  reg rva_in_reg_rw_sva_4;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_4;
  wire GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  wire GBCore_DecodeAxiRead_switch_lp_nor_tmp_1;
  wire GBCore_DecodeAxiRead_switch_lp_equal_tmp_5;
  wire GBCore_DecodeAxiRead_switch_lp_equal_tmp_4;
  wire [2:0] GBCore_PushOutputs_switch_lp_asn_itm_1_mx0;
  reg rva_in_reg_rw_sva_st_4;
  reg [2:0] GBCore_PushOutputs_switch_lp_asn_itm_3;
  reg while_stage_0_5;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  reg GBCore_DecodeAxiRead_switch_lp_nor_13_itm_2;
  reg GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_2;
  reg GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_1;
  reg while_stage_0_4;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1;
  reg while_stage_0_6;
  reg rva_in_reg_rw_sva_st_3;
  reg rva_in_reg_rw_sva_3;
  reg GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
  reg GBCore_DecodeAxiRead_switch_lp_nor_13_itm_3;
  reg rva_in_reg_rw_sva_st_2;
  reg GBCore_PushOutputs_switch_lp_equal_tmp_1;
  reg [2:0] GBCore_PushOutputs_switch_lp_asn_itm_1;
  reg rva_in_reg_rw_sva_1;
  reg GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
  reg GBCore_DecodeAxiRead_switch_lp_nor_13_itm_1;
  reg [2:0] GBCore_PushOutputs_switch_lp_asn_itm_4;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_15_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_16_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_14_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_15_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_13_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_14_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_12_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_13_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_12_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_11_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_11_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_10_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_10_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_9_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_9_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_8_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_8_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_7_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_6_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_5_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_4_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_3_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_2_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_1;
  reg large_mem_write_arbxbar_xbar_for_1_1_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_4_itm_1;
  reg large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_1;
  reg while_stage_0_7;
  reg while_and_11_itm_1;
  reg crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  reg while_stage_0_3;
  wire large_mem_banks_write_if_for_if_mux_cse;
  wire large_mem_banks_write_if_for_if_mux_1_cse;
  wire large_mem_banks_read_for_mux_cse;
  wire large_mem_banks_read_for_mux_1_cse;
  wire large_mem_banks_write_if_for_if_mux_4_cse;
  wire large_mem_banks_write_if_for_if_mux_5_cse;
  wire large_mem_banks_read_for_mux_4_cse;
  wire large_mem_banks_read_for_mux_5_cse;
  wire large_mem_banks_write_if_for_if_mux_8_cse;
  wire large_mem_banks_write_if_for_if_mux_9_cse;
  wire large_mem_banks_read_for_mux_8_cse;
  wire large_mem_banks_read_for_mux_9_cse;
  wire large_mem_banks_write_if_for_if_mux_12_cse;
  wire large_mem_banks_write_if_for_if_mux_13_cse;
  wire large_mem_banks_read_for_mux_12_cse;
  wire large_mem_banks_read_for_mux_13_cse;
  wire large_mem_banks_write_if_for_if_mux_16_cse;
  wire large_mem_banks_write_if_for_if_mux_17_cse;
  wire large_mem_banks_read_for_mux_16_cse;
  wire large_mem_banks_read_for_mux_17_cse;
  wire large_mem_banks_write_if_for_if_mux_20_cse;
  wire large_mem_banks_write_if_for_if_mux_21_cse;
  wire large_mem_banks_read_for_mux_20_cse;
  wire large_mem_banks_read_for_mux_21_cse;
  wire large_mem_banks_write_if_for_if_mux_24_cse;
  wire large_mem_banks_write_if_for_if_mux_25_cse;
  wire large_mem_banks_read_for_mux_24_cse;
  wire large_mem_banks_read_for_mux_25_cse;
  wire large_mem_banks_write_if_for_if_mux_28_cse;
  wire large_mem_banks_write_if_for_if_mux_29_cse;
  wire large_mem_banks_read_for_mux_28_cse;
  wire large_mem_banks_read_for_mux_29_cse;
  wire large_mem_banks_write_if_for_if_mux_32_cse;
  wire large_mem_banks_write_if_for_if_mux_33_cse;
  wire large_mem_banks_read_for_mux_32_cse;
  wire large_mem_banks_read_for_mux_33_cse;
  wire large_mem_banks_write_if_for_if_mux_36_cse;
  wire large_mem_banks_write_if_for_if_mux_37_cse;
  wire large_mem_banks_read_for_mux_36_cse;
  wire large_mem_banks_read_for_mux_37_cse;
  wire large_mem_banks_write_if_for_if_mux_40_cse;
  wire large_mem_banks_write_if_for_if_mux_41_cse;
  wire large_mem_banks_read_for_mux_40_cse;
  wire large_mem_banks_read_for_mux_41_cse;
  wire large_mem_banks_write_if_for_if_mux_44_cse;
  wire large_mem_banks_write_if_for_if_mux_45_cse;
  wire large_mem_banks_read_for_mux_44_cse;
  wire large_mem_banks_read_for_mux_45_cse;
  wire large_mem_banks_write_if_for_if_mux_48_cse;
  wire large_mem_banks_write_if_for_if_mux_49_cse;
  wire large_mem_banks_read_for_mux_48_cse;
  wire large_mem_banks_read_for_mux_49_cse;
  wire large_mem_banks_write_if_for_if_mux_52_cse;
  wire large_mem_banks_write_if_for_if_mux_53_cse;
  wire large_mem_banks_read_for_mux_52_cse;
  wire large_mem_banks_read_for_mux_53_cse;
  wire large_mem_banks_write_if_for_if_mux_56_cse;
  wire large_mem_banks_write_if_for_if_mux_57_cse;
  wire large_mem_banks_read_for_mux_56_cse;
  wire large_mem_banks_read_for_mux_57_cse;
  wire large_mem_banks_write_if_for_if_mux_60_cse;
  wire large_mem_banks_write_if_for_if_mux_61_cse;
  wire large_mem_banks_read_for_mux_60_cse;
  wire large_mem_banks_read_for_mux_61_cse;
  reg reg_large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_nmp_large_rsp_Push_mioi_iswt0_cse;
  reg reg_rva_out_large_Push_mioi_iswt0_cse;
  reg reg_nmp_large_req_PopNB_mioi_iswt0_cse;
  reg reg_rva_in_large_PopNB_mioi_iswt0_cse;
  wire rva_out_reg_data_and_1_cse;
  wire base_large_and_cse;
  wire and_195_cse;
  wire and_192_cse;
  wire and_189_cse;
  wire and_186_cse;
  wire and_183_cse;
  wire and_180_cse;
  wire and_177_cse;
  wire and_174_cse;
  wire and_171_cse;
  wire and_168_cse;
  wire and_165_cse;
  wire and_162_cse;
  wire and_159_cse;
  wire and_156_cse;
  wire and_153_cse;
  wire and_150_cse;
  wire GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse;
  wire mux_7_tmp;
  wire base_large_or_cse;
  wire GBCore_DecodeAxiRead_switch_lp_or_4_cse;
  wire GBCore_DecodeAxiRead_switch_lp_and_6_cse;
  wire GBCore_DecodeAxiRead_switch_lp_and_7_cse;
  wire GBCore_DecodeAxiRead_switch_lp_and_8_cse;
  wire and_143_rmff;
  wire and_140_rmff;
  wire and_137_rmff;
  wire and_134_rmff;
  wire and_131_rmff;
  wire and_128_rmff;
  wire and_125_rmff;
  wire and_122_rmff;
  wire and_119_rmff;
  wire and_116_rmff;
  wire and_113_rmff;
  wire and_110_rmff;
  wire and_107_rmff;
  wire and_104_rmff;
  wire and_101_rmff;
  wire and_98_rmff;
  wire and_147_rmff;
  wire and_146_rmff;
  wire and_145_rmff;
  reg [7:0] rva_out_reg_data_1_127_120_sva_dfm_3_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000;
  reg [7:0] rva_out_reg_data_1_119_112_sva_dfm_3_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000;
  reg [7:0] rva_out_reg_data_1_103_96_sva_dfm_3_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000000;
  reg [7:0] rva_out_reg_data_1_95_88_sva_dfm_3_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000000;
  reg [7:0] rva_out_reg_data_1_87_80_sva_dfm_3_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000000;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000000;
  reg [7:0] rva_out_reg_data_1_71_64_sva_dfm_3_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000000;
  reg [7:0] rva_out_reg_data_1_63_56_sva_dfm_3_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000000;
  reg [7:0] rva_out_reg_data_1_55_48_sva_dfm_3_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000000;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000000;
  reg [7:0] rva_out_reg_data_1_39_32_sva_dfm_3_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000000;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000000;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000000;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi000000;
  reg [7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_7_0;
  wire [7:0] rva_out_reg_data_1_31_0_sva_dfm_1_15_8_1;
  reg [7:0] rva_out_reg_data_1_31_0_sva_dfm_3_7_0;
  wire [7:0] rva_out_reg_data_1_31_0_sva_dfm_1_7_0_1;
  reg [7:0] large_port_read_out_data_0_0_sva_dfm_1;
  reg [7:0] large_req_reg_vector_index_sva_1_1;
  reg [15:0] large_req_reg_timestep_index_sva_1;
  reg [7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_7_0;
  reg [7:0] large_write_data_data_0_15_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_14_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_13_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_12_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_11_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_10_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_9_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_8_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_7_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_6_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_5_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_4_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_3_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_2_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_1_lpi_1_dfm_4_2_16;
  reg [7:0] large_write_data_data_0_0_lpi_1_dfm_4_2_16;
  wire [15:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_1_mx0w1;
  reg [15:0] while_if_while_if_and_1_itm_3;
  wire [15:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_2_mx0w1;
  reg [15:0] while_if_while_if_and_3_itm_3;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi_1;
  reg [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112_lpi_1;
  reg [7:0] large_port_read_out_data_0_0_sva;
  reg [7:0] num_vector_large_1_sva;
  reg [7:0] num_vector_large_2_sva;
  reg [7:0] num_vector_large_3_sva;
  reg [15:0] base_large_1_sva;
  reg [15:0] base_large_2_sva;
  reg GBCore_DecodeAxiWrite_switch_lp_equal_tmp_2;
  reg GBCore_DecodeAxiRead_switch_lp_equal_tmp_3;
  reg [7:0] rva_out_reg_data_1_55_48_sva_dfm_1_1;
  reg [7:0] rva_out_reg_data_1_55_48_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_1_55_48_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_1_55_48_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_1_63_56_sva_dfm_1_1;
  reg [7:0] rva_out_reg_data_1_63_56_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_1_63_56_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_1_63_56_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_1_87_80_sva_dfm_1_1;
  reg [7:0] rva_out_reg_data_1_87_80_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_1_87_80_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_1_87_80_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_1_95_88_sva_dfm_1_1;
  reg [7:0] rva_out_reg_data_1_95_88_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_1_95_88_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_1_95_88_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_1_119_112_sva_dfm_1_1;
  reg [7:0] rva_out_reg_data_1_119_112_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_1_119_112_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_1_119_112_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_1_127_120_sva_dfm_1_1;
  reg [7:0] rva_out_reg_data_1_127_120_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_1_127_120_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_1_127_120_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_1_39_32_sva_dfm_1_1;
  reg [7:0] rva_out_reg_data_1_39_32_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_1_39_32_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_1_39_32_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_1_71_64_sva_dfm_1_1;
  reg [7:0] rva_out_reg_data_1_71_64_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_1_71_64_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_1_71_64_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_1_103_96_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_1_103_96_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_1_103_96_sva_dfm_1_4;
  reg GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
  reg GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
  reg large_req_reg_is_write_sva_1;
  reg large_req_reg_is_write_sva_2;
  reg [15:0] GBCore_SetLargeBuffer_1U_base_addr_acc_3_1;
  reg large_read_req_valid_0_lpi_1_dfm_3_1;
  reg large_read_req_valid_0_lpi_1_dfm_3_2;
  reg [7:0] large_write_data_data_0_0_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_1_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_2_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_3_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_4_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_5_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_6_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_7_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_8_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_9_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_10_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_11_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_12_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_13_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_14_lpi_1_dfm_4_1;
  reg [7:0] large_write_data_data_0_15_lpi_1_dfm_4_1;
  reg [7:0] num_vector_large_0_sva_dfm_3_1;
  reg [7:0] num_vector_large_1_sva_dfm_3_1;
  reg [7:0] num_vector_large_2_sva_dfm_3_1;
  reg [7:0] num_vector_large_3_sva_dfm_3_1;
  reg [15:0] base_large_0_sva_dfm_3_1;
  reg [15:0] base_large_1_sva_dfm_3_1;
  reg [15:0] base_large_2_sva_dfm_3_1;
  reg [15:0] large_mem_write_arbxbar_xbar_for_empty_sva_1;
  reg [3:0] crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1;
  reg GBCore_PushOutputs_switch_lp_equal_tmp_2;
  reg GBCore_DecodeAxiRead_switch_lp_nor_13_itm_4;
  reg GBCore_DecodeAxiRead_switch_lp_nor_13_itm_5;
  reg [2:0] while_if_while_if_and_itm_1;
  reg [15:0] while_if_while_if_and_1_itm_2;
  reg [15:0] while_if_while_if_and_3_itm_2;
  reg [7:0] while_if_while_if_and_5_itm_1;
  reg [7:0] while_if_while_if_and_6_itm_1;
  reg [7:0] while_if_while_if_and_7_itm_1;
  reg [7:0] while_if_while_if_and_8_itm_1;
  reg [7:0] while_if_while_if_and_9_itm_1;
  reg [7:0] while_if_while_if_and_10_itm_1;
  reg [7:0] while_if_while_if_and_11_itm_1;
  reg [7:0] while_if_while_if_and_12_itm_1;
  reg [7:0] while_if_while_if_and_13_itm_1;
  reg [7:0] while_if_while_if_and_14_itm_1;
  reg [7:0] while_if_while_if_and_15_itm_1;
  reg [7:0] while_if_while_if_and_16_itm_1;
  reg [7:0] while_if_while_if_and_17_itm_1;
  reg [7:0] while_if_while_if_and_18_itm_1;
  reg [7:0] while_if_while_if_and_19_itm_1;
  reg [7:0] while_if_while_if_and_20_itm_1;
  reg while_mux_11_itm_1;
  reg while_mux_11_itm_2;
  reg GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_2;
  reg [2:0] GBCore_PushOutputs_switch_lp_asn_itm_2;
  reg [15:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_31_16;
  reg [7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_7_0;
  reg [7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_3_7_0;
  reg [7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_7_0;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi_1_mx0;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000002;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000002;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000002;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000002;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000002;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000002;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000002;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000002;
  wire [7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000002;
  wire [7:0] large_port_read_out_data_0_0_sva_mx0;
  wire [7:0] num_vector_large_0_sva_mx0;
  wire [7:0] num_vector_large_1_sva_mx1;
  wire [7:0] num_vector_large_2_sva_mx1;
  wire [7:0] num_vector_large_3_sva_mx1;
  wire [15:0] base_large_0_sva_mx0;
  wire [15:0] base_large_1_sva_mx1;
  wire [15:0] base_large_2_sva_mx1;
  wire [2:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_mx0w1;
  wire [15:0] GBCore_SetLargeBuffer_1U_base_addr_sva_1;
  wire [16:0] nl_GBCore_SetLargeBuffer_1U_base_addr_sva_1;
  wire [15:0] large_write_addrs_lpi_1_dfm_6;
  wire [3:0] large_read_addrs_0_lpi_1_dfm_4_mx1_3_0;
  wire base_large_and_3_ssc;
  reg [7:0] base_large_3_sva_15_8;
  reg [7:0] base_large_3_sva_7_0;
  reg [7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_24;
  reg [7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_23_16;
  wire [7:0] base_large_3_sva_mx2_15_8;
  wire [7:0] base_large_3_sva_mx2_7_0;
  reg [7:0] reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_0;
  reg [7:0] reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_1;
  wire GBCore_SetLargeBuffer_1U_base_addr_and_ssc;
  wire GBCore_DecodeAxiRead_switch_lp_and_16_ssc;
  reg [7:0] reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_31_16_ftd;
  reg [7:0] reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_31_16_ftd_1;
  reg [7:0] base_large_3_sva_dfm_3_1_15_8;
  reg [7:0] base_large_3_sva_dfm_3_1_7_0;
  reg [7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_31_24;
  reg [7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_23_16;
  wire GBCore_DecodeAxiRead_switch_lp_and_13_cse;
  wire rva_out_reg_data_and_10_cse;
  wire GBCore_PushOutputs_switch_lp_and_cse;
  wire large_mem_write_arbxbar_xbar_for_1_for_and_cse;
  wire large_req_reg_is_write_and_cse;
  wire large_write_data_data_and_cse;
  wire while_if_and_cse;
  wire large_req_reg_vector_index_and_cse;
  wire GBCore_DecodeAxiRead_switch_lp_and_15_cse;
  wire large_mem_write_arbxbar_xbar_for_empty_and_cse;
  wire while_if_and_3_cse;
  wire while_if_and_6_cse;
  wire while_if_and_4_cse;
  wire while_if_and_8_cse;
  wire rva_out_reg_data_and_19_cse;
  wire GBCore_DecodeAxiRead_switch_lp_and_21_cse;
  wire rva_out_reg_data_and_28_cse;
  wire GBCore_DecodeAxiRead_switch_lp_and_25_cse;
  wire GBCore_DecodeAxiRead_switch_lp_and_23_cse;
  wire [7:0] rva_out_reg_data_1_31_0_sva_dfm_1_31_24;
  wire [7:0] rva_out_reg_data_1_31_0_sva_dfm_1_23_16;
  wire data_in_tmp_operator_for_and_32_cse;
  wire data_in_tmp_operator_for_and_33_cse;
  wire and_214_cse;
  wire and_223_cse;
  wire and_286_cse;
  wire and_334_cse;
  wire and_363_cse;
  wire and_549_cse;
  wire nand_17_cse;
  wire and_cse;
  reg reg_rva_out_reg_data_1_127_120_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_1_119_112_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_1_103_96_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_1_95_88_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_1_39_32_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_1_87_80_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_1_55_48_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_1_71_64_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_1_63_56_sva_dfm_1_4_enexo;
  reg reg_large_write_data_data_0_15_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_14_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_13_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_12_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_11_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_10_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_9_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_8_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_7_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_6_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_5_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_4_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_3_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_2_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_1_lpi_1_dfm_4_1_enexo;
  reg reg_large_write_data_data_0_0_lpi_1_dfm_4_1_enexo;
  reg reg_while_if_while_if_and_3_itm_2_enexo;
  reg reg_while_if_while_if_and_1_itm_2_enexo;
  reg reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_enexo;
  reg reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_1_enexo;
  reg reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_3_7_0_enexo;
  reg reg_base_large_2_enexo;
  reg reg_base_large_1_enexo;
  reg reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_7_0_enexo;
  reg reg_rva_out_reg_data_1_103_96_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_1_71_64_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_1_39_32_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_1_127_120_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_1_119_112_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_1_95_88_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_1_87_80_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_1_63_56_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_1_55_48_sva_dfm_1_2_enexo;
  reg reg_base_large_3_1_enexo;
  reg reg_rva_out_reg_data_1_71_64_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_1_39_32_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_1_127_120_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_1_119_112_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_1_95_88_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_1_87_80_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_1_63_56_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_1_55_48_sva_dfm_1_1_enexo;
  reg reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_16_enexo;
  reg reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_16_1_enexo;
  reg reg_base_large_3_sva_dfm_3_1_enexo;
  wire rva_out_reg_data_and_45_enex5;
  wire rva_out_reg_data_and_46_enex5;
  wire rva_out_reg_data_and_47_enex5;
  wire rva_out_reg_data_and_48_enex5;
  wire rva_out_reg_data_and_49_enex5;
  wire rva_out_reg_data_and_50_enex5;
  wire rva_out_reg_data_and_51_enex5;
  wire rva_out_reg_data_and_52_enex5;
  wire rva_out_reg_data_and_53_enex5;
  wire large_write_data_data_and_32_enex5;
  wire large_write_data_data_and_33_enex5;
  wire large_write_data_data_and_34_enex5;
  wire large_write_data_data_and_35_enex5;
  wire large_write_data_data_and_36_enex5;
  wire large_write_data_data_and_37_enex5;
  wire large_write_data_data_and_38_enex5;
  wire large_write_data_data_and_39_enex5;
  wire large_write_data_data_and_40_enex5;
  wire large_write_data_data_and_41_enex5;
  wire large_write_data_data_and_42_enex5;
  wire large_write_data_data_and_43_enex5;
  wire large_write_data_data_and_44_enex5;
  wire large_write_data_data_and_45_enex5;
  wire large_write_data_data_and_46_enex5;
  wire large_write_data_data_and_47_enex5;
  wire while_if_and_25_enex5;
  wire while_if_and_26_enex5;
  wire GBCore_DecodeAxiRead_switch_lp_and_29_enex5;
  wire GBCore_DecodeAxiRead_switch_lp_and_30_enex5;
  wire GBCore_DecodeAxiRead_switch_lp_and_31_enex5;
  wire while_if_and_27_enex5;
  wire while_if_and_28_enex5;
  wire GBCore_DecodeAxiRead_switch_lp_and_20_enex5;
  wire rva_out_reg_data_and_54_enex5;
  wire rva_out_reg_data_and_55_enex5;
  wire rva_out_reg_data_and_56_enex5;
  wire rva_out_reg_data_and_57_enex5;
  wire rva_out_reg_data_and_58_enex5;
  wire rva_out_reg_data_and_59_enex5;
  wire rva_out_reg_data_and_60_enex5;
  wire rva_out_reg_data_and_61_enex5;
  wire rva_out_reg_data_and_62_enex5;
  wire rva_out_reg_data_and_63_enex5;
  wire rva_out_reg_data_and_64_enex5;
  wire rva_out_reg_data_and_65_enex5;
  wire rva_out_reg_data_and_66_enex5;
  wire rva_out_reg_data_and_67_enex5;
  wire rva_out_reg_data_and_68_enex5;
  wire rva_out_reg_data_and_69_enex5;
  wire rva_out_reg_data_and_70_enex5;
  wire rva_out_reg_data_and_71_enex5;
  wire GBCore_SetLargeBuffer_1U_base_addr_and_2_enex5;
  wire GBCore_SetLargeBuffer_1U_base_addr_and_3_enex5;
  wire base_large_and_8_enex5;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_11;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_13;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_28;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_28;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_28;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_28;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_29;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_29;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_29;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_29;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_30;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_30;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_30;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_30;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_15;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_31;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_31;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_31;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_31;
  wire mux_6_nl;
  wire mux_8_nl;
  wire mux_nl;
  wire nor_6_nl;
  wire nor_7_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_1_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_o000000;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_262_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_16_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_264_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_32_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_266_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_48_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_268_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_64_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_270_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_80_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_272_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_96_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_274_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_112_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_276_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_128_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_278_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_144_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_280_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_160_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_282_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_176_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_284_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_192_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_286_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_208_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_256_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_224_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_258_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_240_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_260_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000000;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_1_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_333_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_17_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_348_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_33_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_363_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_49_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_378_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_65_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_393_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_81_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_408_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_97_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_423_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_113_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_438_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_129_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_453_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_145_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_468_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_161_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_483_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_177_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_498_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_193_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_513_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_209_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_288_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_225_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_303_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_241_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_318_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000001;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_13_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_345_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_29_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_360_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_45_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_375_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_61_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_390_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_77_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_405_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_93_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_420_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_109_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_435_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_125_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_450_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_141_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_465_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_157_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_480_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_173_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_495_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_189_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_510_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_205_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_525_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_221_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_300_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_237_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_315_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_253_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_330_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000002;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_2_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_334_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_18_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_349_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_34_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_364_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_50_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_379_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_66_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_394_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_82_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_409_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_98_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_424_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_114_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_439_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_130_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_454_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_146_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_469_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_162_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_484_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_178_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_499_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_194_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_514_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_210_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_289_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_226_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_304_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_242_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_319_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000003;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_3_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_335_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_19_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_350_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_35_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_365_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_51_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_380_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_67_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_395_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_83_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_410_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_99_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_425_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_115_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_440_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_131_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_455_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_147_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_470_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_163_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_485_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_179_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_500_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_195_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_515_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_211_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_290_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_227_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_305_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_243_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_320_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000004;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_5_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_337_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_21_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_352_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_37_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_367_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_53_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_382_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_69_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_397_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_85_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_412_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_101_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_427_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_117_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_442_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_133_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_457_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_149_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_472_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_165_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_487_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_181_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_502_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_197_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_517_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_213_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_292_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_229_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_307_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_245_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_322_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000005;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_9_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_341_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_25_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_356_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_41_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_371_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_57_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_386_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_73_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_401_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_89_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_416_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_105_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_431_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_121_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_446_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_137_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_461_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_153_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_476_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_169_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_491_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_185_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_506_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_201_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_521_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_217_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_296_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_233_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_311_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_249_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_326_nl;
  wire GBCore_PollNMPPort_GBCore_PollNMPPort_and_20_nl;
  wire while_if_while_if_and_5_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_21_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_22_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_23_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_24_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_25_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_26_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_27_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_28_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_29_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_30_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_31_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_32_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_33_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_34_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_35_nl;
  wire[7:0] GBCore_PollNMPPort_GBCore_PollNMPPort_and_36_nl;
  wire GBCore_PollNMPPort_GBCore_PollNMPPort_nor_1_nl;
  wire while_if_while_if_and_6_nl;
  wire[15:0] while_if_while_if_and_1_nl;
  wire rva_in_reg_rw_not_42_nl;
  wire[15:0] while_if_while_if_and_3_nl;
  wire or_85_nl;
  wire mux_3_nl;
  wire nand_4_nl;
  wire or_nl;
  wire mux_5_nl;
  wire nor_11_nl;
  wire mux_4_nl;
  wire nor_12_nl;
  wire nand_5_nl;
  wire and_209_nl;
  wire mux_9_nl;
  wire nor_100_nl;
  wire[15:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_21_nl;
  wire GBCore_DecodeAxiRead_switch_lp_not_20_nl;
  wire[7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_20_nl;
  wire GBCore_DecodeAxiRead_switch_lp_not_19_nl;
  wire[2:0] GBCore_DecodeAxiRead_switch_lp_mux1h_20_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000006;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_15_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_347_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_31_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_362_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_47_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_377_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_63_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_392_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_79_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_407_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_95_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_422_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_111_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_437_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_127_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_452_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_143_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_467_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_159_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_482_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_175_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_497_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_191_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_512_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_207_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_527_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_223_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_302_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_239_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_317_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_255_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_332_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000007;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_14_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_346_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_30_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_361_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_46_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_376_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_62_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_391_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_78_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_406_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_94_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_421_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_110_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_436_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_126_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_451_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_142_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_466_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_158_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_481_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_174_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_496_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_190_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_511_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_206_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_526_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_222_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_301_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_238_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_316_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_254_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_331_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000008;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_12_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_344_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_28_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_359_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_44_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_374_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_60_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_389_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_76_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_404_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_92_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_419_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_108_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_434_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_124_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_449_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_140_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_464_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_156_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_479_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_172_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_494_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_188_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_509_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_204_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_524_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_220_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_299_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_236_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_314_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_252_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_329_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000009;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_11_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_343_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_27_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_358_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_43_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_373_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_59_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_388_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_75_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_403_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_91_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_418_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_107_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_433_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_123_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_448_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_139_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_463_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_155_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_478_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_171_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_493_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_187_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_508_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_203_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_523_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_219_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_298_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_235_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_313_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_251_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_328_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000010;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_4_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_336_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_20_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_351_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_36_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_366_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_52_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_381_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_68_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_396_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_84_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_411_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_100_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_426_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_116_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_441_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_132_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_456_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_148_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_471_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_164_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_486_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_180_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_501_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_196_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_516_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_212_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_291_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_228_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_306_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_244_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_321_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000011;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_10_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_342_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_26_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_357_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_42_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_372_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_58_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_387_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_74_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_402_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_90_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_417_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_106_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_432_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_122_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_447_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_138_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_462_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_154_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_477_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_170_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_492_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_186_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_507_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_202_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_522_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_218_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_297_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_234_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_312_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_250_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_327_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000012;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_6_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_338_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_22_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_353_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_38_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_368_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_54_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_383_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_70_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_398_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_86_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_413_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_102_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_428_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_118_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_443_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_134_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_458_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_150_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_473_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_166_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_488_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_182_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_503_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_198_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_518_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_214_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_293_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_230_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_308_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_246_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_323_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000013;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_8_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_340_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_24_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_355_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_40_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_370_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_56_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_385_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_72_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_400_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_88_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_415_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_104_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_430_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_120_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_445_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_136_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_460_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_152_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_475_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_168_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_490_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_184_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_505_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_200_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_520_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_216_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_295_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_232_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_310_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_248_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_325_nl;
  wire[7:0] crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000014;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_7_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_339_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_23_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_354_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_39_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_369_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_55_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_384_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_71_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_399_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_87_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_414_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_103_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_429_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_119_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_444_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_135_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_459_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_151_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_474_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_167_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_489_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_183_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_504_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_199_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_519_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_215_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_294_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_231_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_309_nl;
  wire[7:0] large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_247_nl;
  wire large_mem_write_arbxbar_xbar_for_1_for_not_324_nl;
  wire large_req_reg_is_write_not_18_nl;
  wire[7:0] GBCore_DecodeAxiRead_switch_lp_mux_11_nl;
  wire[7:0] GBCore_DecodeAxiRead_switch_lp_mux_12_nl;
  wire[7:0] GBCore_DecodeAxiRead_switch_lp_mux_10_nl;
  wire mux_2_nl;
  wire nor_nl;
  wire mux_1_nl;
  wire nor_14_nl;
  wire nand_6_nl;
  wire and_210_nl;
  wire[7:0] GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_7_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [3:0] nl_large_mem_write_arbxbar_xbar_for_lshift_rg_s;
  assign nl_large_mem_write_arbxbar_xbar_for_lshift_rg_s = MUX_v_4_2_2((GBCore_PollNMPPort_GBCore_PollNMPPort_and_2_mx0w1[3:0]),
      (while_if_while_if_and_3_itm_3[3:0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  wire[7:0] rva_out_reg_data_mux_8_nl;
  wire[7:0] rva_out_reg_data_mux_7_nl;
  wire[7:0] data_in_tmp_operator_for_data_in_tmp_operator_for_and_2_nl;
  wire GBCore_PushOutputs_switch_lp_not_3_nl;
  wire[7:0] rva_out_reg_data_mux_6_nl;
  wire[7:0] rva_out_reg_data_mux_5_nl;
  wire[7:0] rva_out_reg_data_mux_4_nl;
  wire[7:0] data_in_tmp_operator_for_data_in_tmp_operator_for_and_1_nl;
  wire GBCore_PushOutputs_switch_lp_not_2_nl;
  wire[7:0] rva_out_reg_data_mux_3_nl;
  wire[7:0] rva_out_reg_data_mux_2_nl;
  wire[7:0] rva_out_reg_data_mux_1_nl;
  wire[7:0] data_in_tmp_operator_for_data_in_tmp_operator_for_and_nl;
  wire GBCore_PushOutputs_switch_lp_not_nl;
  wire[7:0] rva_out_reg_data_mux_nl;
  wire[7:0] data_in_tmp_operator_for_data_in_tmp_operator_for_mux1h_1_nl;
  wire[7:0] data_in_tmp_operator_for_data_in_tmp_operator_for_mux1h_2_nl;
  wire[7:0] data_in_tmp_operator_for_data_in_tmp_operator_for_mux1h_nl;
  wire[7:0] large_port_read_out_data_large_port_read_out_data_mux1h_nl;
  wire large_port_read_out_data_large_port_read_out_data_nor_nl;
  wire large_port_read_out_data_and_1_nl;
  wire [127:0] nl_GBCore_GBCoreRun_rva_out_large_Push_mioi_inst_rva_out_large_Push_mioi_m_data_rsc_dat_GBCoreRun;
  assign rva_out_reg_data_mux_8_nl = MUX_v_8_2_2(rva_out_reg_data_1_127_120_sva_dfm_3_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000,
      and_dcpl_94);
  assign rva_out_reg_data_mux_7_nl = MUX_v_8_2_2(rva_out_reg_data_1_119_112_sva_dfm_3_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000,
      and_dcpl_94);
  assign GBCore_PushOutputs_switch_lp_not_3_nl = ~ and_dcpl_95;
  assign data_in_tmp_operator_for_data_in_tmp_operator_for_and_2_nl = MUX_v_8_2_2(8'b00000000,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000,
      GBCore_PushOutputs_switch_lp_not_3_nl);
  assign rva_out_reg_data_mux_6_nl = MUX_v_8_2_2(rva_out_reg_data_1_103_96_sva_dfm_3_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000000,
      and_dcpl_94);
  assign rva_out_reg_data_mux_5_nl = MUX_v_8_2_2(rva_out_reg_data_1_95_88_sva_dfm_3_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000000,
      and_dcpl_94);
  assign rva_out_reg_data_mux_4_nl = MUX_v_8_2_2(rva_out_reg_data_1_87_80_sva_dfm_3_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000000,
      and_dcpl_94);
  assign GBCore_PushOutputs_switch_lp_not_2_nl = ~ and_dcpl_95;
  assign data_in_tmp_operator_for_data_in_tmp_operator_for_and_1_nl = MUX_v_8_2_2(8'b00000000,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000000,
      GBCore_PushOutputs_switch_lp_not_2_nl);
  assign rva_out_reg_data_mux_3_nl = MUX_v_8_2_2(rva_out_reg_data_1_71_64_sva_dfm_3_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000000,
      and_dcpl_94);
  assign rva_out_reg_data_mux_2_nl = MUX_v_8_2_2(rva_out_reg_data_1_63_56_sva_dfm_3_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000000,
      and_dcpl_94);
  assign rva_out_reg_data_mux_1_nl = MUX_v_8_2_2(rva_out_reg_data_1_55_48_sva_dfm_3_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000000,
      and_dcpl_94);
  assign GBCore_PushOutputs_switch_lp_not_nl = ~ and_dcpl_95;
  assign data_in_tmp_operator_for_data_in_tmp_operator_for_and_nl = MUX_v_8_2_2(8'b00000000,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000000,
      GBCore_PushOutputs_switch_lp_not_nl);
  assign rva_out_reg_data_mux_nl = MUX_v_8_2_2(rva_out_reg_data_1_39_32_sva_dfm_3_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000000,
      and_dcpl_94);
  assign data_in_tmp_operator_for_data_in_tmp_operator_for_mux1h_1_nl = MUX1HOT_v_8_3_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000000,
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_31_24,
      rva_out_reg_data_1_31_0_sva_dfm_1_31_24, {(~ and_dcpl_93) , data_in_tmp_operator_for_and_32_cse
      , data_in_tmp_operator_for_and_33_cse});
  assign data_in_tmp_operator_for_data_in_tmp_operator_for_mux1h_2_nl = MUX1HOT_v_8_3_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000000,
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_23_16,
      rva_out_reg_data_1_31_0_sva_dfm_1_23_16, {(~ and_dcpl_93) , data_in_tmp_operator_for_and_32_cse
      , data_in_tmp_operator_for_and_33_cse});
  assign data_in_tmp_operator_for_data_in_tmp_operator_for_mux1h_nl = MUX1HOT_v_8_3_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi000000,
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_7_0,
      rva_out_reg_data_1_31_0_sva_dfm_1_15_8_1, {(~ and_dcpl_93) , data_in_tmp_operator_for_and_32_cse
      , data_in_tmp_operator_for_and_33_cse});
  assign large_port_read_out_data_large_port_read_out_data_nor_nl = ~(while_and_11_itm_1
      | mux_7_tmp);
  assign large_port_read_out_data_and_1_nl = while_and_11_itm_1 & (~ mux_7_tmp);
  assign large_port_read_out_data_large_port_read_out_data_mux1h_nl = MUX1HOT_v_8_3_2(rva_out_reg_data_1_31_0_sva_dfm_3_7_0,
      rva_out_reg_data_1_31_0_sva_dfm_1_7_0_1, large_port_read_out_data_0_0_sva_dfm_1,
      {large_port_read_out_data_large_port_read_out_data_nor_nl , large_port_read_out_data_and_1_nl
      , mux_7_tmp});
  assign nl_GBCore_GBCoreRun_rva_out_large_Push_mioi_inst_rva_out_large_Push_mioi_m_data_rsc_dat_GBCoreRun
      = {rva_out_reg_data_mux_8_nl , rva_out_reg_data_mux_7_nl , data_in_tmp_operator_for_data_in_tmp_operator_for_and_2_nl
      , rva_out_reg_data_mux_6_nl , rva_out_reg_data_mux_5_nl , rva_out_reg_data_mux_4_nl
      , data_in_tmp_operator_for_data_in_tmp_operator_for_and_1_nl , rva_out_reg_data_mux_3_nl
      , rva_out_reg_data_mux_2_nl , rva_out_reg_data_mux_1_nl , data_in_tmp_operator_for_data_in_tmp_operator_for_and_nl
      , rva_out_reg_data_mux_nl , data_in_tmp_operator_for_data_in_tmp_operator_for_mux1h_1_nl
      , data_in_tmp_operator_for_data_in_tmp_operator_for_mux1h_2_nl , data_in_tmp_operator_for_data_in_tmp_operator_for_mux1h_nl
      , large_port_read_out_data_large_port_read_out_data_mux1h_nl};
  wire [127:0] nl_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_inst_nmp_large_rsp_Push_mioi_m_read_vector_data_data_rsc_dat_GBCoreRun;
  assign nl_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_inst_nmp_large_rsp_Push_mioi_m_read_vector_data_data_rsc_dat_GBCoreRun
      = {crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000000
      , crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi000000
      , large_port_read_out_data_0_0_sva_dfm_1};
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) large_mem_write_arbxbar_xbar_for_lshift_rg (
      .a(while_mux_11_itm_2),
      .s(nl_large_mem_write_arbxbar_xbar_for_lshift_rg_s[3:0]),
      .z(large_mem_write_arbxbar_xbar_for_lshift_tmp)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd16)) large_mem_read_arbxbar_xbar_for_1_lshift_rg (
      .a(large_read_req_valid_0_lpi_1_dfm_3_2),
      .s(large_read_addrs_0_lpi_1_dfm_4_mx1_3_0),
      .z(large_mem_read_arbxbar_xbar_for_1_lshift_tmp)
    );
  GBModule_GBCore_GBCoreRun_rva_in_large_PopNB_mioi GBCore_GBCoreRun_rva_in_large_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_large_vld(rva_in_large_vld),
      .rva_in_large_rdy(rva_in_large_rdy),
      .rva_in_large_dat(rva_in_large_dat),
      .GBCoreRun_wen(GBCoreRun_wen),
      .GBCoreRun_wten(GBCoreRun_wten),
      .rva_in_large_PopNB_mioi_oswt(reg_rva_in_large_PopNB_mioi_iswt0_cse),
      .rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_large_PopNB_mioi_return_rsc_z_mxwt(rva_in_large_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_large_PopNB_mioi_oswt_pff(fsm_output)
    );
  GBModule_GBCore_GBCoreRun_nmp_large_req_PopNB_mioi GBCore_GBCoreRun_nmp_large_req_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .nmp_large_req_vld(nmp_large_req_vld),
      .nmp_large_req_rdy(nmp_large_req_rdy),
      .nmp_large_req_dat(nmp_large_req_dat),
      .GBCoreRun_wen(GBCoreRun_wen),
      .GBCoreRun_wten(GBCoreRun_wten),
      .nmp_large_req_PopNB_mioi_oswt(reg_nmp_large_req_PopNB_mioi_iswt0_cse),
      .nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt(nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_return_rsc_z_mxwt(nmp_large_req_PopNB_mioi_return_rsc_z_mxwt),
      .nmp_large_req_PopNB_mioi_oswt_pff(and_147_rmff)
    );
  GBModule_GBCore_GBCoreRun_rva_out_large_Push_mioi GBCore_GBCoreRun_rva_out_large_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_large_vld(rva_out_large_vld),
      .rva_out_large_rdy(rva_out_large_rdy),
      .rva_out_large_dat(rva_out_large_dat),
      .GBCoreRun_wen(GBCoreRun_wen),
      .rva_out_large_Push_mioi_oswt(reg_rva_out_large_Push_mioi_iswt0_cse),
      .rva_out_large_Push_mioi_wen_comp(rva_out_large_Push_mioi_wen_comp),
      .rva_out_large_Push_mioi_m_data_rsc_dat_GBCoreRun(nl_GBCore_GBCoreRun_rva_out_large_Push_mioi_inst_rva_out_large_Push_mioi_m_data_rsc_dat_GBCoreRun[127:0]),
      .rva_out_large_Push_mioi_oswt_pff(and_146_rmff)
    );
  GBModule_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .nmp_large_rsp_vld(nmp_large_rsp_vld),
      .nmp_large_rsp_rdy(nmp_large_rsp_rdy),
      .nmp_large_rsp_dat(nmp_large_rsp_dat),
      .GBCoreRun_wen(GBCoreRun_wen),
      .nmp_large_rsp_Push_mioi_oswt(reg_nmp_large_rsp_Push_mioi_iswt0_cse),
      .nmp_large_rsp_Push_mioi_wen_comp(nmp_large_rsp_Push_mioi_wen_comp),
      .nmp_large_rsp_Push_mioi_m_read_vector_data_data_rsc_dat_GBCoreRun(nl_GBCore_GBCoreRun_nmp_large_rsp_Push_mioi_inst_nmp_large_rsp_Push_mioi_m_read_vector_data_data_rsc_dat_GBCoreRun[127:0]),
      .nmp_large_rsp_Push_mioi_oswt_pff(and_145_rmff)
    );
  GBModule_GBCore_GBCoreRun_wait_dp GBCore_GBCoreRun_wait_dp_inst (
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d),
      .GBCoreRun_wen(GBCoreRun_wen),
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo(reg_large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo_ir_unreg(and_143_rmff),
      .large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo(reg_large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo_ir_unreg(and_140_rmff),
      .large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo(reg_large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo_ir_unreg(and_137_rmff),
      .large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo(reg_large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo_ir_unreg(and_134_rmff),
      .large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo(reg_large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo_ir_unreg(and_131_rmff),
      .large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo(reg_large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo_ir_unreg(and_128_rmff),
      .large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo(reg_large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo_ir_unreg(and_125_rmff),
      .large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo(reg_large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo_ir_unreg(and_122_rmff),
      .large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo(reg_large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo_ir_unreg(and_119_rmff),
      .large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo(reg_large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo_ir_unreg(and_116_rmff),
      .large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo(reg_large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo_ir_unreg(and_113_rmff),
      .large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo(reg_large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo_ir_unreg(and_110_rmff),
      .large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo(reg_large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo_ir_unreg(and_107_rmff),
      .large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo(reg_large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo_ir_unreg(and_104_rmff),
      .large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo(reg_large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo_ir_unreg(and_101_rmff),
      .large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo(reg_large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo_ir_cse),
      .large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo_ir_unreg(and_98_rmff)
    );
  GBModule_GBCore_GBCoreRun_staller GBCore_GBCoreRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .GBCoreRun_wen(GBCoreRun_wen),
      .GBCoreRun_wten(GBCoreRun_wten),
      .rva_out_large_Push_mioi_wen_comp(rva_out_large_Push_mioi_wen_comp),
      .nmp_large_rsp_Push_mioi_wen_comp(nmp_large_rsp_Push_mioi_wen_comp)
    );
  GBModule_GBCore_GBCoreRun_GBCoreRun_fsm GBCore_GBCoreRun_GBCoreRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .GBCoreRun_wen(GBCoreRun_wen),
      .fsm_output(fsm_output)
    );
  assign large_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_195_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = large_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl large_mem_banks_load_store_for_1_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign large_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_195_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = large_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = large_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_1_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = large_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = large_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_1_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = large_mem_banks_write_if_for_if_mux_1_cse;
  assign large_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_24);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = large_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_1_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign large_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_24);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = large_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = large_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_1_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = large_mem_banks_read_for_mux_1_cse;
  assign large_mem_banks_write_if_for_if_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_192_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 = large_mem_banks_write_if_for_if_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_2_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 );
  assign large_mem_banks_write_if_for_if_mux_5_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_192_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2 = large_mem_banks_write_if_for_if_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 = large_mem_banks_write_if_for_if_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_2_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2 = large_mem_banks_write_if_for_if_mux_5_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1
      = large_mem_banks_write_if_for_if_mux_4_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_2_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1
      = large_mem_banks_write_if_for_if_mux_5_cse;
  assign large_mem_banks_read_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_26);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 = large_mem_banks_read_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_2_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 );
  assign large_mem_banks_read_for_mux_5_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_26);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3 = large_mem_banks_read_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 = large_mem_banks_read_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_2_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3 = large_mem_banks_read_for_mux_5_cse;
  assign large_mem_banks_write_if_for_if_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_189_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 = large_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_3_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 );
  assign large_mem_banks_write_if_for_if_mux_9_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_189_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4 = large_mem_banks_write_if_for_if_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 = large_mem_banks_write_if_for_if_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_3_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4 = large_mem_banks_write_if_for_if_mux_9_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2
      = large_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_3_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2
      = large_mem_banks_write_if_for_if_mux_9_cse;
  assign large_mem_banks_read_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_28);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 = large_mem_banks_read_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_3_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 );
  assign large_mem_banks_read_for_mux_9_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_28);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5 = large_mem_banks_read_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 = large_mem_banks_read_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_3_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5 = large_mem_banks_read_for_mux_9_cse;
  assign large_mem_banks_write_if_for_if_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_186_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 = large_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_4_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 );
  assign large_mem_banks_write_if_for_if_mux_13_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_186_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6 = large_mem_banks_write_if_for_if_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 = large_mem_banks_write_if_for_if_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_4_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6 = large_mem_banks_write_if_for_if_mux_13_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3
      = large_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_4_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3
      = large_mem_banks_write_if_for_if_mux_13_cse;
  assign large_mem_banks_read_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_30);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 = large_mem_banks_read_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_4_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 );
  assign large_mem_banks_read_for_mux_13_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_30);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7 = large_mem_banks_read_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 = large_mem_banks_read_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_4_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7 = large_mem_banks_read_for_mux_13_cse;
  assign large_mem_banks_write_if_for_if_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_183_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 = large_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_5_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 );
  assign large_mem_banks_write_if_for_if_mux_17_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_183_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8 = large_mem_banks_write_if_for_if_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 = large_mem_banks_write_if_for_if_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_5_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8 = large_mem_banks_write_if_for_if_mux_17_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4
      = large_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_5_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4
      = large_mem_banks_write_if_for_if_mux_17_cse;
  assign large_mem_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_32);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 = large_mem_banks_read_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_5_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 );
  assign large_mem_banks_read_for_mux_17_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_32);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9 = large_mem_banks_read_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 = large_mem_banks_read_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_5_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9 = large_mem_banks_read_for_mux_17_cse;
  assign large_mem_banks_write_if_for_if_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_180_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 = large_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_6_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 );
  assign large_mem_banks_write_if_for_if_mux_21_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_180_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10 = large_mem_banks_write_if_for_if_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 = large_mem_banks_write_if_for_if_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_6_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10 = large_mem_banks_write_if_for_if_mux_21_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5
      = large_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_6_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5
      = large_mem_banks_write_if_for_if_mux_21_cse;
  assign large_mem_banks_read_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_34);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 = large_mem_banks_read_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_6_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 );
  assign large_mem_banks_read_for_mux_21_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_34);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11 = large_mem_banks_read_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 = large_mem_banks_read_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_6_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11 = large_mem_banks_read_for_mux_21_cse;
  assign large_mem_banks_write_if_for_if_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_177_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 = large_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_7_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 );
  assign large_mem_banks_write_if_for_if_mux_25_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_177_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12 = large_mem_banks_write_if_for_if_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 = large_mem_banks_write_if_for_if_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_7_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12 = large_mem_banks_write_if_for_if_mux_25_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6
      = large_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_7_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6
      = large_mem_banks_write_if_for_if_mux_25_cse;
  assign large_mem_banks_read_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_36);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 = large_mem_banks_read_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_7_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 );
  assign large_mem_banks_read_for_mux_25_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_36);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13 = large_mem_banks_read_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 = large_mem_banks_read_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_7_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13 = large_mem_banks_read_for_mux_25_cse;
  assign large_mem_banks_write_if_for_if_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_174_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 = large_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_8_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 );
  assign large_mem_banks_write_if_for_if_mux_29_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_174_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14 = large_mem_banks_write_if_for_if_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 = large_mem_banks_write_if_for_if_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_8_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14 = large_mem_banks_write_if_for_if_mux_29_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7
      = large_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_8_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7
      = large_mem_banks_write_if_for_if_mux_29_cse;
  assign large_mem_banks_read_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_38);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 = large_mem_banks_read_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_8_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 );
  assign large_mem_banks_read_for_mux_29_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_38);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15 = large_mem_banks_read_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 = large_mem_banks_read_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_8_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15 = large_mem_banks_read_for_mux_29_cse;
  assign large_mem_banks_write_if_for_if_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, and_171_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 = large_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_9_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 );
  assign large_mem_banks_write_if_for_if_mux_33_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_171_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16 = large_mem_banks_write_if_for_if_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 = large_mem_banks_write_if_for_if_mux_32_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_9_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16 = large_mem_banks_write_if_for_if_mux_33_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8
      = large_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_9_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8
      = large_mem_banks_write_if_for_if_mux_33_cse;
  assign large_mem_banks_read_for_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_40);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 = large_mem_banks_read_for_mux_32_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_9_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 );
  assign large_mem_banks_read_for_mux_33_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_40);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17 = large_mem_banks_read_for_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 = large_mem_banks_read_for_mux_32_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_9_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17 = large_mem_banks_read_for_mux_33_cse;
  assign large_mem_banks_write_if_for_if_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, and_168_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 = large_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_10_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 );
  assign large_mem_banks_write_if_for_if_mux_37_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_168_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18 = large_mem_banks_write_if_for_if_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 = large_mem_banks_write_if_for_if_mux_36_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_10_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18 = large_mem_banks_write_if_for_if_mux_37_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9
      = large_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_10_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9
      = large_mem_banks_write_if_for_if_mux_37_cse;
  assign large_mem_banks_read_for_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_42);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 = large_mem_banks_read_for_mux_36_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_10_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 );
  assign large_mem_banks_read_for_mux_37_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_42);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19 = large_mem_banks_read_for_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 = large_mem_banks_read_for_mux_36_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_10_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19 = large_mem_banks_read_for_mux_37_cse;
  assign large_mem_banks_write_if_for_if_mux_40_cse = MUX1HOT_s_1_1_2(1'b1, and_165_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 = large_mem_banks_write_if_for_if_mux_40_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_11_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 );
  assign large_mem_banks_write_if_for_if_mux_41_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_165_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20 = large_mem_banks_write_if_for_if_mux_41_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 = large_mem_banks_write_if_for_if_mux_40_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_11_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20 = large_mem_banks_write_if_for_if_mux_41_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_10
      = large_mem_banks_write_if_for_if_mux_40_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_11_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_10  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_10 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_10
      = large_mem_banks_write_if_for_if_mux_41_cse;
  assign large_mem_banks_read_for_mux_40_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_44);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 = large_mem_banks_read_for_mux_40_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_11_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 );
  assign large_mem_banks_read_for_mux_41_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_44);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21 = large_mem_banks_read_for_mux_41_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 = large_mem_banks_read_for_mux_40_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_11_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21 = large_mem_banks_read_for_mux_41_cse;
  assign large_mem_banks_write_if_for_if_mux_44_cse = MUX1HOT_s_1_1_2(1'b1, and_162_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 = large_mem_banks_write_if_for_if_mux_44_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_12_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 );
  assign large_mem_banks_write_if_for_if_mux_45_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_162_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22 = large_mem_banks_write_if_for_if_mux_45_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 = large_mem_banks_write_if_for_if_mux_44_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_12_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22 = large_mem_banks_write_if_for_if_mux_45_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_11
      = large_mem_banks_write_if_for_if_mux_44_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_12_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_11  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_11 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_11
      = large_mem_banks_write_if_for_if_mux_45_cse;
  assign large_mem_banks_read_for_mux_44_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_46);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 = large_mem_banks_read_for_mux_44_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_12_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 );
  assign large_mem_banks_read_for_mux_45_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_46);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23 = large_mem_banks_read_for_mux_45_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 = large_mem_banks_read_for_mux_44_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_12_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23 = large_mem_banks_read_for_mux_45_cse;
  assign large_mem_banks_write_if_for_if_mux_48_cse = MUX1HOT_s_1_1_2(1'b1, and_159_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 = large_mem_banks_write_if_for_if_mux_48_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_13_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 );
  assign large_mem_banks_write_if_for_if_mux_49_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_159_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24 = large_mem_banks_write_if_for_if_mux_49_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 = large_mem_banks_write_if_for_if_mux_48_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_13_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24 = large_mem_banks_write_if_for_if_mux_49_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_12
      = large_mem_banks_write_if_for_if_mux_48_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_13_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_12  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_12 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_12
      = large_mem_banks_write_if_for_if_mux_49_cse;
  assign large_mem_banks_read_for_mux_48_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_48);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 = large_mem_banks_read_for_mux_48_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_13_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 );
  assign large_mem_banks_read_for_mux_49_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_48);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25 = large_mem_banks_read_for_mux_49_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 = large_mem_banks_read_for_mux_48_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_13_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25 = large_mem_banks_read_for_mux_49_cse;
  assign large_mem_banks_write_if_for_if_mux_52_cse = MUX1HOT_s_1_1_2(1'b1, and_156_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 = large_mem_banks_write_if_for_if_mux_52_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_14_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 );
  assign large_mem_banks_write_if_for_if_mux_53_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_156_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26 = large_mem_banks_write_if_for_if_mux_53_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 = large_mem_banks_write_if_for_if_mux_52_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_14_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26 = large_mem_banks_write_if_for_if_mux_53_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_13
      = large_mem_banks_write_if_for_if_mux_52_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_14_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_13  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_13 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_13
      = large_mem_banks_write_if_for_if_mux_53_cse;
  assign large_mem_banks_read_for_mux_52_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_50);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 = large_mem_banks_read_for_mux_52_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_14_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 );
  assign large_mem_banks_read_for_mux_53_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_50);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27 = large_mem_banks_read_for_mux_53_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 = large_mem_banks_read_for_mux_52_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_14_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27 = large_mem_banks_read_for_mux_53_cse;
  assign large_mem_banks_write_if_for_if_mux_56_cse = MUX1HOT_s_1_1_2(1'b1, and_153_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_28 = large_mem_banks_write_if_for_if_mux_56_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_15_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_28  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_28 );
  assign large_mem_banks_write_if_for_if_mux_57_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_153_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_28 = large_mem_banks_write_if_for_if_mux_57_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_28 = large_mem_banks_write_if_for_if_mux_56_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_15_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_28  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_28 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_28 = large_mem_banks_write_if_for_if_mux_57_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_14
      = large_mem_banks_write_if_for_if_mux_56_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_15_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_14  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_14 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_14
      = large_mem_banks_write_if_for_if_mux_57_cse;
  assign large_mem_banks_read_for_mux_56_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_52);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_29 = large_mem_banks_read_for_mux_56_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_15_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_29  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_29 );
  assign large_mem_banks_read_for_mux_57_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_52);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_29 = large_mem_banks_read_for_mux_57_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_29 = large_mem_banks_read_for_mux_56_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_15_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_29  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_29 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_29 = large_mem_banks_read_for_mux_57_cse;
  assign large_mem_banks_write_if_for_if_mux_60_cse = MUX1HOT_s_1_1_2(1'b1, and_150_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_30 = large_mem_banks_write_if_for_if_mux_60_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl large_mem_banks_load_store_for_16_GBCore_GBCoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_30  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_30 );
  assign large_mem_banks_write_if_for_if_mux_61_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen,
      and_150_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_30 = large_mem_banks_write_if_for_if_mux_61_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_30 = large_mem_banks_write_if_for_if_mux_60_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl large_mem_banks_load_store_for_16_GBCore_GBCoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_30  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_30 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_30 = large_mem_banks_write_if_for_if_mux_61_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_15
      = large_mem_banks_write_if_for_if_mux_60_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl large_mem_banks_load_store_for_16_GBCore_GBCoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_15  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_15 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_15
      = large_mem_banks_write_if_for_if_mux_61_cse;
  assign large_mem_banks_read_for_mux_60_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_54);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_31 = large_mem_banks_read_for_mux_60_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl large_mem_banks_load_store_for_16_GBCore_GBCoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_31  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_31 );
  assign large_mem_banks_read_for_mux_61_cse = MUX1HOT_s_1_1_2(GBCoreRun_wen, and_dcpl_54);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_31 = large_mem_banks_read_for_mux_61_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_31 = large_mem_banks_read_for_mux_60_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl large_mem_banks_load_store_for_16_GBCore_GBCoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_31  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_31 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_31 = large_mem_banks_read_for_mux_61_cse;
  assign mux_6_nl = MUX_s_1_2_2((~ (GBCore_PushOutputs_switch_lp_asn_itm_4[2])),
      (GBCore_PushOutputs_switch_lp_asn_itm_4[2]), GBCore_PushOutputs_switch_lp_asn_itm_4[0]);
  assign mux_7_tmp = MUX_s_1_2_2(or_tmp_11, mux_6_nl, fsm_output);
  assign and_98_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[15]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[15]))
      & while_stage_0_5) | ((large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_15_1_itm_1
      | large_mem_write_arbxbar_xbar_for_1_16_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_101_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[14]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[14]))
      & while_stage_0_5) | ((large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_14_1_itm_1
      | large_mem_write_arbxbar_xbar_for_1_15_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_104_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[13]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[13]))
      & while_stage_0_5) | ((large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_13_1_itm_1
      | large_mem_write_arbxbar_xbar_for_1_14_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_107_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[12]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[12]))
      & while_stage_0_5) | ((large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_12_1_itm_1
      | large_mem_write_arbxbar_xbar_for_1_13_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_110_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[11]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[11]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_12_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_11_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_113_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[10]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_11_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_10_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_116_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[9]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[9]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_10_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_9_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_119_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[8]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[8]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_9_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_8_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_122_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[7]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_8_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_125_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[6]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_7_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_128_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[5]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_6_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_131_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[4]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_5_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_134_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[3]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_4_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_137_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[2]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_3_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_140_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[1]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_2_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_143_rmff = ((((large_mem_write_arbxbar_xbar_for_lshift_tmp[0]) | (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]))
      & while_stage_0_5) | ((large_mem_write_arbxbar_xbar_for_1_1_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_4_itm_1
      | large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_1)
      & while_stage_0_6)) & fsm_output;
  assign and_145_rmff = and_dcpl_94 & (GBCore_PushOutputs_switch_lp_asn_itm_4[1])
      & while_stage_0_7;
  assign mux_8_nl = MUX_s_1_2_2((GBCore_PushOutputs_switch_lp_asn_itm_4[2]), (~ or_tmp_11),
      GBCore_PushOutputs_switch_lp_asn_itm_4[1]);
  assign and_146_rmff = mux_8_nl & while_stage_0_7;
  assign and_147_rmff = reg_rva_in_large_PopNB_mioi_iswt0_cse & (~ rva_in_large_PopNB_mioi_return_rsc_z_mxwt);
  assign and_214_cse = ((while_stage_0_7 & while_and_11_itm_1 & (~(GBCore_DecodeAxiRead_switch_lp_nor_13_itm_5
      & GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_5))) | ((~ rva_in_reg_rw_sva_4)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_4
      & while_stage_0_6)) & GBCoreRun_wen;
  assign GBCore_DecodeAxiRead_switch_lp_and_13_cse = GBCoreRun_wen & and_dcpl_1 &
      (~(rva_in_reg_rw_sva_4 | rva_in_reg_rw_sva_st_4));
  assign nor_6_nl = ~((~ (GBCore_PushOutputs_switch_lp_asn_itm_3[2])) | (GBCore_PushOutputs_switch_lp_asn_itm_3[0]));
  assign nor_7_nl = ~((GBCore_PushOutputs_switch_lp_asn_itm_3[2]) | (~ (GBCore_PushOutputs_switch_lp_asn_itm_3[0])));
  assign mux_nl = MUX_s_1_2_2(nor_6_nl, nor_7_nl, GBCore_PushOutputs_switch_lp_asn_itm_3[1]);
  assign rva_out_reg_data_and_10_cse = GBCoreRun_wen & mux_nl & while_stage_0_6;
  assign rva_out_reg_data_and_45_enex5 = rva_out_reg_data_and_10_cse & reg_rva_out_reg_data_1_127_120_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_46_enex5 = rva_out_reg_data_and_10_cse & reg_rva_out_reg_data_1_119_112_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_47_enex5 = rva_out_reg_data_and_10_cse & reg_rva_out_reg_data_1_103_96_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_48_enex5 = rva_out_reg_data_and_10_cse & reg_rva_out_reg_data_1_95_88_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_49_enex5 = rva_out_reg_data_and_10_cse & reg_rva_out_reg_data_1_39_32_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_50_enex5 = rva_out_reg_data_and_10_cse & reg_rva_out_reg_data_1_87_80_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_51_enex5 = rva_out_reg_data_and_10_cse & reg_rva_out_reg_data_1_55_48_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_52_enex5 = rva_out_reg_data_and_10_cse & reg_rva_out_reg_data_1_71_64_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_53_enex5 = rva_out_reg_data_and_10_cse & reg_rva_out_reg_data_1_63_56_sva_dfm_1_4_enexo;
  assign and_223_cse = (((GBCore_PushOutputs_switch_lp_asn_itm_3[0]) & (GBCore_PushOutputs_switch_lp_asn_itm_3[2]))
      | or_dcpl_1) & GBCoreRun_wen & (crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1
      | (~ while_stage_0_7)) & while_stage_0_6;
  assign GBCore_PushOutputs_switch_lp_and_cse = GBCoreRun_wen & while_stage_0_6;
  assign large_mem_write_arbxbar_xbar_for_1_for_and_cse = GBCoreRun_wen & while_stage_0_5;
  assign large_req_reg_is_write_and_cse = GBCoreRun_wen & and_dcpl_55 & GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_1;
  assign large_write_data_data_and_cse = GBCoreRun_wen & while_stage_0_4;
  assign large_write_data_data_and_32_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_15_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_33_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_14_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_34_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_13_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_35_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_12_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_36_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_11_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_37_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_10_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_38_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_9_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_39_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_8_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_40_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_7_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_41_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_6_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_42_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_5_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_43_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_4_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_44_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_3_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_45_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_2_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_46_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_1_lpi_1_dfm_4_1_enexo;
  assign large_write_data_data_and_47_enex5 = large_write_data_data_and_cse & reg_large_write_data_data_0_0_lpi_1_dfm_4_1_enexo;
  assign while_if_and_cse = GBCoreRun_wen & and_dcpl_58;
  assign while_if_and_25_enex5 = while_if_and_cse & reg_while_if_while_if_and_3_itm_2_enexo;
  assign while_if_and_26_enex5 = while_if_and_cse & reg_while_if_while_if_and_1_itm_2_enexo;
  assign large_req_reg_vector_index_and_cse = GBCoreRun_wen & and_dcpl_59 & nmp_large_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_if_and_3_cse = GBCoreRun_wen & while_stage_0_3;
  assign while_if_and_4_cse = GBCoreRun_wen & reg_rva_in_large_PopNB_mioi_iswt0_cse;
  assign and_286_cse = GBCoreRun_wen & or_dcpl_1 & (~ while_stage_0_6) & while_stage_0_7;
  assign GBCore_DecodeAxiRead_switch_lp_and_15_cse = GBCoreRun_wen & and_dcpl_63
      & (~(rva_in_reg_rw_sva_3 | rva_in_reg_rw_sva_st_3));
  assign GBCore_DecodeAxiRead_switch_lp_and_16_ssc = GBCoreRun_wen & and_dcpl_63
      & (~ rva_in_reg_rw_sva_3) & (~ rva_in_reg_rw_sva_st_3) & GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_3
      & GBCore_DecodeAxiRead_switch_lp_nor_13_itm_3;
  assign GBCore_DecodeAxiRead_switch_lp_and_29_enex5 = GBCore_DecodeAxiRead_switch_lp_and_16_ssc
      & reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_enexo;
  assign GBCore_DecodeAxiRead_switch_lp_and_30_enex5 = GBCore_DecodeAxiRead_switch_lp_and_16_ssc
      & reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_1_enexo;
  assign GBCore_DecodeAxiRead_switch_lp_and_31_enex5 = GBCore_DecodeAxiRead_switch_lp_and_16_ssc
      & reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_3_7_0_enexo;
  assign large_mem_write_arbxbar_xbar_for_empty_and_cse = GBCoreRun_wen & while_stage_0_5
      & large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_and_tmp
      & (~ crossbar_spec_GB_Large_WordType_16U_16U_for_mux_tmp);
  assign rva_out_reg_data_and_1_cse = GBCoreRun_wen & ((and_dcpl_63 & (~ rva_in_reg_rw_sva_3))
      | and_dcpl_204);
  assign nand_17_cse = ~(rva_in_large_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_large_PopNB_mioi_iswt0_cse);
  assign and_334_cse = nand_17_cse & fsm_output & while_if_and_3_cse;
  assign while_if_and_6_cse = GBCoreRun_wen & and_dcpl_72;
  assign while_if_and_27_enex5 = while_if_and_6_cse & reg_base_large_2_enexo;
  assign while_if_and_28_enex5 = while_if_and_6_cse & reg_base_large_1_enexo;
  assign base_large_or_cse = and_dcpl_206 | and_cse;
  assign base_large_and_cse = GBCoreRun_wen & base_large_or_cse;
  assign and_363_cse = (~((~((rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[15:0]==16'b0000000000000001)
      & rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt & rva_in_large_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100))) & while_stage_0_3))
      & while_if_and_4_cse;
  assign while_if_and_8_cse = GBCoreRun_wen & and_cse;
  assign GBCore_DecodeAxiRead_switch_lp_and_20_enex5 = GBCoreRun_wen & and_dcpl_58
      & (~ rva_in_reg_rw_sva_st_2) & GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_2
      & GBCore_DecodeAxiRead_switch_lp_nor_13_itm_2 & reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_7_0_enexo;
  assign nand_4_nl = ~((GBCore_PushOutputs_switch_lp_asn_itm_1[1:0]==2'b11));
  assign or_nl = (GBCore_PushOutputs_switch_lp_asn_itm_1[1:0]!=2'b00);
  assign mux_3_nl = MUX_s_1_2_2(nand_4_nl, or_nl, GBCore_PushOutputs_switch_lp_asn_itm_1[2]);
  assign rva_out_reg_data_and_19_cse = GBCoreRun_wen & (~(mux_3_nl & GBCore_PushOutputs_switch_lp_equal_tmp_1))
      & and_dcpl_58 & (~ rva_in_reg_rw_sva_st_2);
  assign rva_out_reg_data_and_54_enex5 = rva_out_reg_data_and_19_cse & reg_rva_out_reg_data_1_103_96_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_55_enex5 = rva_out_reg_data_and_19_cse & reg_rva_out_reg_data_1_71_64_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_56_enex5 = rva_out_reg_data_and_19_cse & reg_rva_out_reg_data_1_39_32_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_57_enex5 = rva_out_reg_data_and_19_cse & reg_rva_out_reg_data_1_127_120_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_58_enex5 = rva_out_reg_data_and_19_cse & reg_rva_out_reg_data_1_119_112_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_59_enex5 = rva_out_reg_data_and_19_cse & reg_rva_out_reg_data_1_95_88_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_60_enex5 = rva_out_reg_data_and_19_cse & reg_rva_out_reg_data_1_87_80_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_61_enex5 = rva_out_reg_data_and_19_cse & reg_rva_out_reg_data_1_63_56_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_62_enex5 = rva_out_reg_data_and_19_cse & reg_rva_out_reg_data_1_55_48_sva_dfm_1_2_enexo;
  assign GBCore_DecodeAxiRead_switch_lp_and_21_cse = GBCoreRun_wen & and_dcpl_72
      & (~ rva_in_reg_rw_sva_1);
  assign GBCore_DecodeAxiRead_switch_lp_or_4_cse = (~((nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt!=2'b00)))
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1;
  assign GBCore_DecodeAxiRead_switch_lp_and_6_cse = (nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt==2'b01)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
  assign GBCore_DecodeAxiRead_switch_lp_and_7_cse = (nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt==2'b10)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
  assign GBCore_DecodeAxiRead_switch_lp_and_8_cse = (nmp_large_req_PopNB_mioi_data_memory_index_rsc_z_mxwt==2'b11)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
  assign nor_11_nl = ~((~ nmp_large_req_PopNB_mioi_return_rsc_z_mxwt) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
  assign nor_12_nl = ~(rva_in_reg_rw_sva_1 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1));
  assign nand_5_nl = ~(rva_in_reg_rw_sva_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
  assign mux_4_nl = MUX_s_1_2_2(nor_12_nl, nand_5_nl, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt);
  assign and_209_nl = GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_1 & GBCore_DecodeAxiRead_switch_lp_nor_13_itm_1;
  assign mux_5_nl = MUX_s_1_2_2(nor_11_nl, mux_4_nl, and_209_nl);
  assign GBCore_DecodeAxiRead_switch_lp_and_23_cse = GBCoreRun_wen & mux_5_nl & while_stage_0_3;
  assign rva_out_reg_data_and_28_cse = GBCoreRun_wen & ((while_mux_2_tmp!=3'b101))
      & and_dcpl_72 & (~ rva_in_reg_rw_sva_1);
  assign rva_out_reg_data_and_63_enex5 = rva_out_reg_data_and_28_cse & reg_base_large_3_1_enexo;
  assign rva_out_reg_data_and_64_enex5 = rva_out_reg_data_and_28_cse & reg_rva_out_reg_data_1_71_64_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_65_enex5 = rva_out_reg_data_and_28_cse & reg_rva_out_reg_data_1_39_32_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_66_enex5 = rva_out_reg_data_and_28_cse & reg_rva_out_reg_data_1_127_120_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_67_enex5 = rva_out_reg_data_and_28_cse & reg_rva_out_reg_data_1_119_112_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_68_enex5 = rva_out_reg_data_and_28_cse & reg_rva_out_reg_data_1_95_88_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_69_enex5 = rva_out_reg_data_and_28_cse & reg_rva_out_reg_data_1_87_80_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_70_enex5 = rva_out_reg_data_and_28_cse & reg_rva_out_reg_data_1_63_56_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_71_enex5 = rva_out_reg_data_and_28_cse & reg_rva_out_reg_data_1_55_48_sva_dfm_1_1_enexo;
  assign GBCore_DecodeAxiRead_switch_lp_and_25_cse = GBCoreRun_wen & and_cse & (~
      rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_cse = reg_rva_in_large_PopNB_mioi_iswt0_cse & rva_in_large_PopNB_mioi_return_rsc_z_mxwt;
  assign nor_100_nl = ~((~((rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[15:0]!=16'b0000000000000001)
      | while_stage_0_3)) | (rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]!=4'b0100)
      | rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign mux_9_nl = MUX_s_1_2_2(while_stage_0_3, nor_100_nl, and_cse);
  assign and_549_cse = mux_9_nl & fsm_output & GBCoreRun_wen;
  assign and_150_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[15]);
  assign and_153_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[14]);
  assign and_156_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[13]);
  assign and_159_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[12]);
  assign and_162_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[11]);
  assign and_165_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[10]);
  assign and_168_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[9]);
  assign and_171_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[8]);
  assign and_174_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[7]);
  assign and_177_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[6]);
  assign and_180_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[5]);
  assign and_183_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[4]);
  assign and_186_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[3]);
  assign and_189_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[2]);
  assign and_192_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[1]);
  assign and_195_cse = while_stage_0_5 & (large_mem_write_arbxbar_xbar_for_lshift_tmp[0]);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_347_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_15_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_347_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_362_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_31_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_362_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_377_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_47_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_377_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_392_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_63_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_392_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_407_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_79_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_407_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_422_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_95_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_422_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_437_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_111_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_437_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_452_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_127_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_452_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_467_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_143_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_467_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_482_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_159_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_482_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_497_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_175_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_497_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_512_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_191_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_512_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_527_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_207_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_527_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_302_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_223_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_302_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_317_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_239_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_317_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_332_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_255_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[127:120]),
      large_mem_write_arbxbar_xbar_for_1_for_not_332_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000006
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_15_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_31_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_47_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_63_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_79_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_95_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_111_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_127_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_143_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_159_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_175_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_191_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_207_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_223_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_239_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_255_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000002,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000006,
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_346_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_14_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_346_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_361_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_30_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_361_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_376_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_46_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_376_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_391_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_62_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_391_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_406_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_78_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_406_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_421_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_94_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_421_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_436_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_110_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_436_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_451_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_126_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_451_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_466_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_142_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_466_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_481_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_158_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_481_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_496_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_174_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_496_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_511_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_190_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_511_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_526_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_206_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_526_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_301_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_222_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_301_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_316_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_238_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_316_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_331_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_254_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[119:112]),
      large_mem_write_arbxbar_xbar_for_1_for_not_331_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000007
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_14_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_30_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_46_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_62_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_78_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_94_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_110_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_126_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_142_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_158_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_174_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_190_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_206_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_222_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_238_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_254_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000002,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000007,
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_344_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_12_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_344_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_359_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_28_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_359_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_374_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_44_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_374_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_389_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_60_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_389_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_404_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_76_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_404_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_419_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_92_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_419_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_434_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_108_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_434_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_449_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_124_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_449_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_464_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_140_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_464_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_479_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_156_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_479_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_494_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_172_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_494_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_509_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_188_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_509_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_524_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_204_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_524_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_299_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_220_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_299_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_314_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_236_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_314_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_329_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_252_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[103:96]),
      large_mem_write_arbxbar_xbar_for_1_for_not_329_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000008
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_12_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_28_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_44_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_60_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_76_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_92_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_108_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_124_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_140_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_156_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_172_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_188_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_204_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_220_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_236_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_252_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000002,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000008,
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_343_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_11_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_343_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_358_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_27_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_358_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_373_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_43_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_373_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_388_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_59_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_388_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_403_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_75_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_403_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_418_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_91_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_418_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_433_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_107_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_433_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_448_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_123_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_448_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_463_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_139_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_463_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_478_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_155_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_478_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_493_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_171_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_493_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_508_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_187_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_508_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_523_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_203_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_523_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_298_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_219_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_298_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_313_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_235_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_313_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_328_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_251_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[95:88]),
      large_mem_write_arbxbar_xbar_for_1_for_not_328_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000009
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_11_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_27_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_43_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_59_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_75_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_91_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_107_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_123_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_139_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_155_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_171_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_187_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_203_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_219_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_235_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_251_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000002,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000009,
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_336_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_4_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_336_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_351_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_20_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_351_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_366_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_36_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_366_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_381_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_52_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_381_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_396_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_68_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_396_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_411_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_84_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_411_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_426_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_100_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_426_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_441_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_116_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_441_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_456_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_132_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_456_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_471_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_148_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_471_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_486_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_164_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_486_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_501_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_180_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_501_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_516_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_196_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_516_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_291_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_212_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_291_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_306_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_228_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_306_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_321_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_244_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[39:32]),
      large_mem_write_arbxbar_xbar_for_1_for_not_321_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000010
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_4_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_20_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_36_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_52_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_68_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_84_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_100_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_116_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_132_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_148_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_164_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_180_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_196_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_212_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_228_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_244_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000002,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000010,
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_342_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_10_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_342_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_357_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_26_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_357_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_372_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_42_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_372_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_387_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_58_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_387_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_402_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_74_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_402_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_417_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_90_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_417_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_432_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_106_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_432_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_447_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_122_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_447_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_462_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_138_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_462_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_477_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_154_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_477_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_492_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_170_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_492_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_507_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_186_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_507_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_522_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_202_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_522_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_297_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_218_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_297_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_312_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_234_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_312_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_327_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_250_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[87:80]),
      large_mem_write_arbxbar_xbar_for_1_for_not_327_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000011
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_10_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_26_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_42_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_58_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_74_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_90_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_106_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_122_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_138_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_154_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_170_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_186_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_202_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_218_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_234_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_250_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000002,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000011,
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_338_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_6_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_338_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_353_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_22_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_353_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_368_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_38_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_368_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_383_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_54_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_383_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_398_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_70_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_398_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_413_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_86_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_413_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_428_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_102_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_428_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_443_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_118_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_443_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_458_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_134_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_458_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_473_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_150_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_473_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_488_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_166_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_488_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_503_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_182_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_503_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_518_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_198_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_518_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_293_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_214_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_293_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_308_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_230_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_308_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_323_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_246_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[55:48]),
      large_mem_write_arbxbar_xbar_for_1_for_not_323_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000012
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_6_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_22_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_38_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_54_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_70_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_86_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_102_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_118_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_134_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_150_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_166_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_182_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_198_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_214_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_230_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_246_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000002,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000012,
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_340_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_8_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_340_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_355_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_24_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_355_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_370_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_40_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_370_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_385_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_56_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_385_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_400_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_72_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_400_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_415_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_88_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_415_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_430_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_104_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_430_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_445_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_120_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_445_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_460_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_136_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_460_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_475_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_152_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_475_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_490_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_168_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_490_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_505_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_184_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_505_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_520_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_200_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_520_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_295_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_216_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_295_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_310_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_232_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_310_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_325_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_248_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[71:64]),
      large_mem_write_arbxbar_xbar_for_1_for_not_325_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000013
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_8_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_24_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_40_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_56_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_72_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_88_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_104_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_120_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_136_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_152_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_168_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_184_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_200_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_216_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_232_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_248_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000002,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000013,
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_339_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_7_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_339_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_354_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_23_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_354_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_369_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_39_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_369_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_384_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_55_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_384_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_399_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_71_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_399_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_414_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_87_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_414_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_429_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_103_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_429_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_444_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_119_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_444_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_459_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_135_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_459_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_474_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_151_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_474_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_489_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_167_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_489_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_504_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_183_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_504_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_519_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_199_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_519_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_294_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_215_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_294_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_309_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_231_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_309_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_324_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_247_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[63:56]),
      large_mem_write_arbxbar_xbar_for_1_for_not_324_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000014
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_7_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_23_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_39_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_55_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_71_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_87_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_103_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_119_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_135_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_151_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_167_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_183_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_199_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_215_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_231_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_247_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000002,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000014,
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi_1_mx0
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000002
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000002
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000002
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000002
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000002
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000002
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000002
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000002
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000,
      while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000002
      = MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112_lpi_1,
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000,
      while_stage_0_7);
  assign large_port_read_out_data_0_0_sva_mx0 = MUX_v_8_2_2(large_port_read_out_data_0_0_sva,
      large_port_read_out_data_0_0_sva_dfm_1, while_stage_0_7);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_mux_tmp = MUX_s_1_16_2((large_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (large_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (large_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (large_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[7]), (large_mem_write_arbxbar_xbar_for_lshift_tmp[8]),
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[9]), (large_mem_write_arbxbar_xbar_for_lshift_tmp[10]),
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[11]), (large_mem_write_arbxbar_xbar_for_lshift_tmp[12]),
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[13]), (large_mem_write_arbxbar_xbar_for_lshift_tmp[14]),
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[15]), large_read_addrs_0_lpi_1_dfm_4_mx1_3_0);
  assign num_vector_large_0_sva_mx0 = MUX_v_8_2_2(GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_7_0,
      num_vector_large_0_sva_dfm_3_1, while_stage_0_3);
  assign num_vector_large_1_sva_mx1 = MUX_v_8_2_2(num_vector_large_1_sva, num_vector_large_1_sva_dfm_3_1,
      while_stage_0_3);
  assign num_vector_large_2_sva_mx1 = MUX_v_8_2_2(num_vector_large_2_sva, num_vector_large_2_sva_dfm_3_1,
      while_stage_0_3);
  assign num_vector_large_3_sva_mx1 = MUX_v_8_2_2(num_vector_large_3_sva, num_vector_large_3_sva_dfm_3_1,
      while_stage_0_3);
  assign base_large_0_sva_mx0 = MUX_v_16_2_2(GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_31_16,
      base_large_0_sva_dfm_3_1, while_stage_0_3);
  assign base_large_1_sva_mx1 = MUX_v_16_2_2(base_large_1_sva, base_large_1_sva_dfm_3_1,
      while_stage_0_3);
  assign base_large_2_sva_mx1 = MUX_v_16_2_2(base_large_2_sva, base_large_2_sva_dfm_3_1,
      while_stage_0_3);
  assign GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 = (rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0101);
  assign large_req_reg_is_write_not_18_nl = ~ nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt;
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_mx0w1 = MUX_v_3_2_2(3'b000, ({{2{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}},
      nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}), large_req_reg_is_write_not_18_nl);
  assign GBCore_PushOutputs_switch_lp_asn_itm_1_mx0 = MUX_v_3_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_mx0w1,
      while_if_while_if_and_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
  assign GBCore_DecodeAxiRead_switch_lp_equal_tmp_4 = (rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100);
  assign GBCore_DecodeAxiRead_switch_lp_mux_11_nl = MUX_v_8_2_2((SC_SRAM_CONFIG[31:24]),
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_31_24,
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_5);
  assign rva_out_reg_data_1_31_0_sva_dfm_1_31_24 = MUX_v_8_2_2(8'b00000000, GBCore_DecodeAxiRead_switch_lp_mux_11_nl,
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_5);
  assign GBCore_DecodeAxiRead_switch_lp_mux_12_nl = MUX_v_8_2_2((SC_SRAM_CONFIG[23:16]),
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_23_16,
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_5);
  assign rva_out_reg_data_1_31_0_sva_dfm_1_23_16 = MUX_v_8_2_2(8'b00000000, GBCore_DecodeAxiRead_switch_lp_mux_12_nl,
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_5);
  assign GBCore_DecodeAxiRead_switch_lp_mux_10_nl = MUX_v_8_2_2((SC_SRAM_CONFIG[7:0]),
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_7_0,
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_5);
  assign rva_out_reg_data_1_31_0_sva_dfm_1_7_0_1 = MUX_v_8_2_2(8'b00000000, GBCore_DecodeAxiRead_switch_lp_mux_10_nl,
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_5);
  assign rva_out_reg_data_1_31_0_sva_dfm_1_15_8_1 = (SC_SRAM_CONFIG[15:8]) & (signext_8_1(~
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_5)) & ({{7{GBCore_DecodeAxiRead_switch_lp_nor_13_itm_5}},
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_5});
  assign nl_GBCore_SetLargeBuffer_1U_base_addr_sva_1 = ({reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_0
      , reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_1}) + GBCore_SetLargeBuffer_1U_base_addr_acc_3_1;
  assign GBCore_SetLargeBuffer_1U_base_addr_sva_1 = nl_GBCore_SetLargeBuffer_1U_base_addr_sva_1[15:0];
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_2_mx0w1 = GBCore_SetLargeBuffer_1U_base_addr_sva_1
      & ({{15{large_req_reg_is_write_sva_2}}, large_req_reg_is_write_sva_2}) & ({{15{GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_2}},
      GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_2});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_1_mx0w1 = GBCore_SetLargeBuffer_1U_base_addr_sva_1
      & (signext_16_1(~ large_req_reg_is_write_sva_2)) & ({{15{GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_2}},
      GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_2});
  assign large_read_addrs_0_lpi_1_dfm_4_mx1_3_0 = MUX_v_4_2_2((GBCore_PollNMPPort_GBCore_PollNMPPort_and_1_mx0w1[3:0]),
      (while_if_while_if_and_1_itm_3[3:0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_and_tmp
      = large_read_req_valid_0_lpi_1_dfm_3_2 & ((large_mem_read_arbxbar_xbar_for_1_lshift_tmp!=16'b0000000000000000))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[0]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[0])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[1]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[1])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[2]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[2])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[3]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[3])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[4]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[4])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[5]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[5])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[6]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[6])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[7]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[7])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[8]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[8])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[9]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[9])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[10]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[10])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[11]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[11])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[12]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[12])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[13]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[13])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[14]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[14])))
      & (~((large_mem_write_arbxbar_xbar_for_lshift_tmp[15]) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[15])));
  assign large_write_addrs_lpi_1_dfm_6 = MUX_v_16_2_2(16'b0000000000000000, (rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[15:0]),
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign GBCore_DecodeAxiRead_switch_lp_nor_tmp_1 = ~(GBCore_DecodeAxiRead_switch_lp_equal_tmp_5
      | GBCore_DecodeAxiRead_switch_lp_equal_tmp_4 | GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign GBCore_DecodeAxiRead_switch_lp_equal_tmp_5 = (rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0011);
  assign GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse =
      ~((rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[15:0]==16'b0000000000000001));
  assign while_mux_2_tmp = MUX_v_3_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_mx0w1,
      while_if_while_if_and_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
  assign and_dcpl_1 = while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_4;
  assign or_dcpl_1 = (~(while_stage_0_5 & large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_and_tmp))
      | crossbar_spec_GB_Large_WordType_16U_16U_for_mux_tmp;
  assign and_dcpl_7 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[0]));
  assign and_dcpl_8 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[1]));
  assign and_dcpl_9 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[2]));
  assign and_dcpl_10 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[3]));
  assign and_dcpl_11 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[4]));
  assign and_dcpl_12 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[5]));
  assign and_dcpl_13 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[6]));
  assign and_dcpl_14 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[7]));
  assign and_dcpl_15 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[8]));
  assign and_dcpl_16 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[9]));
  assign and_dcpl_17 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[10]));
  assign and_dcpl_18 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[11]));
  assign and_dcpl_19 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[12]));
  assign and_dcpl_20 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[13]));
  assign and_dcpl_21 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[14]));
  assign and_dcpl_22 = while_stage_0_5 & (~ (large_mem_write_arbxbar_xbar_for_lshift_tmp[15]));
  assign and_dcpl_24 = and_dcpl_7 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign and_dcpl_26 = and_dcpl_8 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign and_dcpl_28 = and_dcpl_9 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign and_dcpl_30 = and_dcpl_10 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign and_dcpl_32 = and_dcpl_11 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign and_dcpl_34 = and_dcpl_12 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign and_dcpl_36 = and_dcpl_13 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign and_dcpl_38 = and_dcpl_14 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign and_dcpl_40 = and_dcpl_15 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[8]);
  assign and_dcpl_42 = and_dcpl_16 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[9]);
  assign and_dcpl_44 = and_dcpl_17 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]);
  assign and_dcpl_46 = and_dcpl_18 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[11]);
  assign and_dcpl_48 = and_dcpl_19 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[12]);
  assign and_dcpl_50 = and_dcpl_20 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[13]);
  assign and_dcpl_52 = and_dcpl_21 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[14]);
  assign and_dcpl_54 = and_dcpl_22 & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[15]);
  assign and_dcpl_55 = while_stage_0_4 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign and_dcpl_58 = while_stage_0_4 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign and_dcpl_59 = while_stage_0_3 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
  assign and_dcpl_63 = while_stage_0_5 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign and_dcpl_72 = while_stage_0_3 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1;
  assign or_tmp_11 = (~ (GBCore_PushOutputs_switch_lp_asn_itm_4[0])) | (GBCore_PushOutputs_switch_lp_asn_itm_4[2]);
  assign and_dcpl_93 = ((GBCore_PushOutputs_switch_lp_asn_itm_4[2]) ^ (GBCore_PushOutputs_switch_lp_asn_itm_4[0]))
      & fsm_output;
  assign and_dcpl_94 = (GBCore_PushOutputs_switch_lp_asn_itm_4[2]) & (GBCore_PushOutputs_switch_lp_asn_itm_4[0]);
  assign and_dcpl_95 = (~((GBCore_PushOutputs_switch_lp_asn_itm_4[2]) & (GBCore_PushOutputs_switch_lp_asn_itm_4[0])))
      & fsm_output;
  assign and_dcpl_199 = ((~(while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_4))
      | rva_in_reg_rw_sva_4) & while_stage_0_7 & while_and_11_itm_1;
  assign and_dcpl_204 = ((~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5)) | rva_in_reg_rw_sva_3) & while_stage_0_6 & GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
  assign and_dcpl_206 = nand_17_cse & while_stage_0_3;
  assign or_dcpl_71 = (rva_in_large_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]!=4'b0100)
      | (~(rva_in_large_PopNB_mioi_return_rsc_z_mxwt & rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt))
      | GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse;
  assign GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_a = GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_7_0;
  assign GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_b = {(large_req_reg_timestep_index_sva_1[15:4])
      , 4'b0000};
  assign GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_c = {large_req_reg_vector_index_sva_1_1
      , (large_req_reg_timestep_index_sva_1[3:0])};
  assign large_mem_banks_bank_a0_a0_a0_a0_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_pff = MUX_v_12_2_2((GBCore_PollNMPPort_GBCore_PollNMPPort_and_1_mx0w1[15:4]),
      (while_if_while_if_and_1_itm_3[15:4]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign large_mem_banks_bank_a0_a0_a0_a0_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[0])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_pff = MUX_v_12_2_2((GBCore_PollNMPPort_GBCore_PollNMPPort_and_2_mx0w1[15:4]),
      (while_if_while_if_and_3_itm_3[15:4]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign large_mem_banks_bank_a0_a0_a0_a0_a_rsci_we_d_pff = and_195_cse;
  assign large_mem_banks_bank_a0_a0_a0_a1_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a0_a0_a0_a1_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[1])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign large_mem_banks_bank_a0_a0_a0_a1_a_rsci_we_d_pff = and_192_cse;
  assign large_mem_banks_bank_a0_a0_a1_a0_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a0_a0_a1_a0_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[2])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign large_mem_banks_bank_a0_a0_a1_a0_a_rsci_we_d_pff = and_189_cse;
  assign large_mem_banks_bank_a0_a0_a1_a1_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a0_a0_a1_a1_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[3])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign large_mem_banks_bank_a0_a0_a1_a1_a_rsci_we_d_pff = and_186_cse;
  assign large_mem_banks_bank_a0_a1_a0_a0_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a0_a1_a0_a0_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[4])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign large_mem_banks_bank_a0_a1_a0_a0_a_rsci_we_d_pff = and_183_cse;
  assign large_mem_banks_bank_a0_a1_a0_a1_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a0_a1_a0_a1_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[5])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign large_mem_banks_bank_a0_a1_a0_a1_a_rsci_we_d_pff = and_180_cse;
  assign large_mem_banks_bank_a0_a1_a1_a0_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a0_a1_a1_a0_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[6])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign large_mem_banks_bank_a0_a1_a1_a0_a_rsci_we_d_pff = and_177_cse;
  assign large_mem_banks_bank_a0_a1_a1_a1_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a0_a1_a1_a1_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[7])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign large_mem_banks_bank_a0_a1_a1_a1_a_rsci_we_d_pff = and_174_cse;
  assign large_mem_banks_bank_a1_a0_a0_a0_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a1_a0_a0_a0_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[8])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[8]);
  assign large_mem_banks_bank_a1_a0_a0_a0_a_rsci_we_d_pff = and_171_cse;
  assign large_mem_banks_bank_a1_a0_a0_a1_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a1_a0_a0_a1_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[9])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[9]);
  assign large_mem_banks_bank_a1_a0_a0_a1_a_rsci_we_d_pff = and_168_cse;
  assign large_mem_banks_bank_a1_a0_a1_a0_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a1_a0_a1_a0_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[10])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[10]);
  assign large_mem_banks_bank_a1_a0_a1_a0_a_rsci_we_d_pff = and_165_cse;
  assign large_mem_banks_bank_a1_a0_a1_a1_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a1_a0_a1_a1_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[11])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[11]);
  assign large_mem_banks_bank_a1_a0_a1_a1_a_rsci_we_d_pff = and_162_cse;
  assign large_mem_banks_bank_a1_a1_a0_a0_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a1_a1_a0_a0_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[12])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[12]);
  assign large_mem_banks_bank_a1_a1_a0_a0_a_rsci_we_d_pff = and_159_cse;
  assign large_mem_banks_bank_a1_a1_a0_a1_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a1_a1_a0_a1_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[13])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[13]);
  assign large_mem_banks_bank_a1_a1_a0_a1_a_rsci_we_d_pff = and_156_cse;
  assign large_mem_banks_bank_a1_a1_a1_a0_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a1_a1_a1_a0_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[14])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[14]);
  assign large_mem_banks_bank_a1_a1_a1_a0_a_rsci_we_d_pff = and_153_cse;
  assign large_mem_banks_bank_a1_a1_a1_a1_a_rsci_d_d = {large_write_data_data_0_15_lpi_1_dfm_4_2_16
      , large_write_data_data_0_14_lpi_1_dfm_4_2_16 , large_write_data_data_0_13_lpi_1_dfm_4_2_16
      , large_write_data_data_0_12_lpi_1_dfm_4_2_16 , large_write_data_data_0_11_lpi_1_dfm_4_2_16
      , large_write_data_data_0_10_lpi_1_dfm_4_2_16 , large_write_data_data_0_9_lpi_1_dfm_4_2_16
      , large_write_data_data_0_8_lpi_1_dfm_4_2_16 , large_write_data_data_0_7_lpi_1_dfm_4_2_16
      , large_write_data_data_0_6_lpi_1_dfm_4_2_16 , large_write_data_data_0_5_lpi_1_dfm_4_2_16
      , large_write_data_data_0_4_lpi_1_dfm_4_2_16 , large_write_data_data_0_3_lpi_1_dfm_4_2_16
      , large_write_data_data_0_2_lpi_1_dfm_4_2_16 , large_write_data_data_0_1_lpi_1_dfm_4_2_16
      , large_write_data_data_0_0_lpi_1_dfm_4_2_16};
  assign large_mem_banks_bank_a1_a1_a1_a1_a_rsci_re_d_pff = while_stage_0_5 & (~
      (large_mem_write_arbxbar_xbar_for_lshift_tmp[15])) & (large_mem_read_arbxbar_xbar_for_1_lshift_tmp[15]);
  assign large_mem_banks_bank_a1_a1_a1_a1_a_rsci_we_d_pff = and_150_cse;
  assign nor_nl = ~((~ GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_1)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign nor_14_nl = ~(rva_in_reg_rw_sva_st_2 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2));
  assign nand_6_nl = ~(rva_in_reg_rw_sva_st_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign mux_1_nl = MUX_s_1_2_2(nor_14_nl, nand_6_nl, GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_1);
  assign and_210_nl = GBCore_DecodeAxiRead_switch_lp_nor_13_itm_2 & GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_2;
  assign mux_2_nl = MUX_s_1_2_2(nor_nl, mux_1_nl, and_210_nl);
  assign GBCore_SetLargeBuffer_1U_base_addr_and_ssc = GBCoreRun_wen & mux_2_nl &
      while_stage_0_4;
  assign GBCore_SetLargeBuffer_1U_base_addr_and_2_enex5 = GBCore_SetLargeBuffer_1U_base_addr_and_ssc
      & reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_16_enexo;
  assign GBCore_SetLargeBuffer_1U_base_addr_and_3_enex5 = GBCore_SetLargeBuffer_1U_base_addr_and_ssc
      & reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_16_1_enexo;
  assign base_large_and_3_ssc = GBCoreRun_wen & base_large_or_cse & fsm_output &
      (nand_17_cse | (~ rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt));
  assign base_large_and_8_enex5 = base_large_and_3_ssc & reg_base_large_3_sva_dfm_3_1_enexo;
  assign base_large_3_sva_mx2_15_8 = MUX_v_8_2_2(base_large_3_sva_15_8, base_large_3_sva_dfm_3_1_15_8,
      while_stage_0_3);
  assign base_large_3_sva_mx2_7_0 = MUX_v_8_2_2(base_large_3_sva_7_0, base_large_3_sva_dfm_3_1_7_0,
      while_stage_0_3);
  assign data_in_tmp_operator_for_and_32_cse = (~ while_and_11_itm_1) & and_dcpl_93;
  assign data_in_tmp_operator_for_and_33_cse = while_and_11_itm_1 & and_dcpl_93;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_nmp_large_rsp_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_out_large_Push_mioi_iswt0_cse <= 1'b0;
      reg_nmp_large_req_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_large_PopNB_mioi_iswt0_cse <= 1'b0;
      while_stage_0_3 <= 1'b0;
      while_stage_0_4 <= 1'b0;
      while_stage_0_5 <= 1'b0;
      while_stage_0_6 <= 1'b0;
      while_stage_0_7 <= 1'b0;
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= 1'b0;
    end
    else if ( GBCoreRun_wen ) begin
      reg_large_mem_banks_bank_a1_a1_a1_a1_a_rsci_cgo_ir_cse <= and_98_rmff;
      reg_large_mem_banks_bank_a1_a1_a1_a0_a_rsci_cgo_ir_cse <= and_101_rmff;
      reg_large_mem_banks_bank_a1_a1_a0_a1_a_rsci_cgo_ir_cse <= and_104_rmff;
      reg_large_mem_banks_bank_a1_a1_a0_a0_a_rsci_cgo_ir_cse <= and_107_rmff;
      reg_large_mem_banks_bank_a1_a0_a1_a1_a_rsci_cgo_ir_cse <= and_110_rmff;
      reg_large_mem_banks_bank_a1_a0_a1_a0_a_rsci_cgo_ir_cse <= and_113_rmff;
      reg_large_mem_banks_bank_a1_a0_a0_a1_a_rsci_cgo_ir_cse <= and_116_rmff;
      reg_large_mem_banks_bank_a1_a0_a0_a0_a_rsci_cgo_ir_cse <= and_119_rmff;
      reg_large_mem_banks_bank_a0_a1_a1_a1_a_rsci_cgo_ir_cse <= and_122_rmff;
      reg_large_mem_banks_bank_a0_a1_a1_a0_a_rsci_cgo_ir_cse <= and_125_rmff;
      reg_large_mem_banks_bank_a0_a1_a0_a1_a_rsci_cgo_ir_cse <= and_128_rmff;
      reg_large_mem_banks_bank_a0_a1_a0_a0_a_rsci_cgo_ir_cse <= and_131_rmff;
      reg_large_mem_banks_bank_a0_a0_a1_a1_a_rsci_cgo_ir_cse <= and_134_rmff;
      reg_large_mem_banks_bank_a0_a0_a1_a0_a_rsci_cgo_ir_cse <= and_137_rmff;
      reg_large_mem_banks_bank_a0_a0_a0_a1_a_rsci_cgo_ir_cse <= and_140_rmff;
      reg_large_mem_banks_bank_a0_a0_a0_a0_a_rsci_cgo_ir_cse <= and_143_rmff;
      reg_nmp_large_rsp_Push_mioi_iswt0_cse <= and_145_rmff;
      reg_rva_out_large_Push_mioi_iswt0_cse <= and_146_rmff;
      reg_nmp_large_req_PopNB_mioi_iswt0_cse <= and_147_rmff;
      reg_rva_in_large_PopNB_mioi_iswt0_cse <= fsm_output;
      while_stage_0_3 <= reg_rva_in_large_PopNB_mioi_iswt0_cse;
      while_stage_0_4 <= while_stage_0_3;
      while_stage_0_5 <= while_stage_0_4;
      while_stage_0_6 <= while_stage_0_5;
      while_stage_0_7 <= while_stage_0_6;
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= MUX_s_1_2_2(GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_2,
          GBCore_PushOutputs_switch_lp_equal_tmp_2, or_85_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_31_24
          <= 8'b00000000;
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_23_16
          <= 8'b00000000;
    end
    else if ( and_214_cse ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_31_24
          <= MUX_v_8_2_2(reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_31_16_ftd,
          rva_out_reg_data_1_31_0_sva_dfm_1_31_24, and_dcpl_199);
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_23_16
          <= MUX_v_8_2_2(reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_31_16_ftd_1,
          rva_out_reg_data_1_31_0_sva_dfm_1_23_16, and_dcpl_199);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= 1'b0;
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_5 <= 1'b0;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_13_cse ) begin
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_5 <= GBCore_DecodeAxiRead_switch_lp_nor_13_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_7_0
          <= 8'b00000000;
    end
    else if ( GBCoreRun_wen & ((and_dcpl_1 & (~ rva_in_reg_rw_sva_4)) | and_dcpl_199)
        ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_5_7_0
          <= MUX_v_8_2_2(GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_7_0,
          rva_out_reg_data_1_31_0_sva_dfm_1_15_8_1, and_dcpl_199);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_127_120_sva_dfm_3_1 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_45_enex5 ) begin
      rva_out_reg_data_1_127_120_sva_dfm_3_1 <= rva_out_reg_data_1_127_120_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_31_0_sva_dfm_3_7_0 <= 8'b00000000;
    end
    else if ( GBCoreRun_wen & while_stage_0_7 & while_and_11_itm_1 ) begin
      rva_out_reg_data_1_31_0_sva_dfm_3_7_0 <= rva_out_reg_data_1_31_0_sva_dfm_1_7_0_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_119_112_sva_dfm_3_1 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_46_enex5 ) begin
      rva_out_reg_data_1_119_112_sva_dfm_3_1 <= rva_out_reg_data_1_119_112_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_103_96_sva_dfm_3_1 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_47_enex5 ) begin
      rva_out_reg_data_1_103_96_sva_dfm_3_1 <= rva_out_reg_data_1_103_96_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_95_88_sva_dfm_3_1 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_48_enex5 ) begin
      rva_out_reg_data_1_95_88_sva_dfm_3_1 <= rva_out_reg_data_1_95_88_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_39_32_sva_dfm_3_1 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_49_enex5 ) begin
      rva_out_reg_data_1_39_32_sva_dfm_3_1 <= rva_out_reg_data_1_39_32_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_87_80_sva_dfm_3_1 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_50_enex5 ) begin
      rva_out_reg_data_1_87_80_sva_dfm_3_1 <= rva_out_reg_data_1_87_80_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_55_48_sva_dfm_3_1 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_51_enex5 ) begin
      rva_out_reg_data_1_55_48_sva_dfm_3_1 <= rva_out_reg_data_1_55_48_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_71_64_sva_dfm_3_1 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_52_enex5 ) begin
      rva_out_reg_data_1_71_64_sva_dfm_3_1 <= rva_out_reg_data_1_71_64_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_63_56_sva_dfm_3_1 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_53_enex5 ) begin
      rva_out_reg_data_1_63_56_sva_dfm_3_1 <= rva_out_reg_data_1_63_56_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000
          <= 8'b00000000;
      large_port_read_out_data_0_0_sva_dfm_1 <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000000
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000000
          <= 8'b00000000;
    end
    else if ( and_223_cse ) begin
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000000
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000001;
      large_port_read_out_data_0_0_sva_dfm_1 <= MUX_v_8_2_2(large_port_read_out_data_0_0_sva_mx0,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_1_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_o000000,
          crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi000000
          <= MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi_1_mx0,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000000,
          crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000
          <= MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000001,
          crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000000
          <= MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000001,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000002,
          crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000000
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000000
          <= MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000001,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000003,
          crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000000
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000000
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000000
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000000
          <= MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000001,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000004,
          crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000000
          <= MUX_v_8_2_2(crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000001,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000005,
          crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1);
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000000
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000000
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000000
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000001;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_PushOutputs_switch_lp_asn_itm_4 <= 3'b000;
      while_and_11_itm_1 <= 1'b0;
    end
    else if ( GBCore_PushOutputs_switch_lp_and_cse ) begin
      GBCore_PushOutputs_switch_lp_asn_itm_4 <= GBCore_PushOutputs_switch_lp_asn_itm_3;
      while_and_11_itm_1 <= (~ rva_in_reg_rw_sva_4) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_7 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_8 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_9 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[2];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_10 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[3];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_11 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[4];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_12 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[5];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_13 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_14 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[7];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_8_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_15 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_8_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[8];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_9_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_16 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_9_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[9];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_10_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_17 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_10_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[10];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_11_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_18 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_11_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[11];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_12_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_19 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_12_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[12];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_13_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_20 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_13_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[13];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_14_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_21 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_14_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[14];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_15_1_itm_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_22 ) begin
      large_mem_read_arbxbar_xbar_requests_transpose_slc_large_mem_read_arbxbar_xbar_requests_transpose_0_15_1_itm_1
          <= large_mem_read_arbxbar_xbar_for_1_lshift_tmp[15];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_write_arbxbar_xbar_for_1_16_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_15_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_14_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_13_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_12_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_11_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_10_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_9_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_8_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_7_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_6_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_5_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_4_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_3_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_2_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= 1'b0;
      large_mem_write_arbxbar_xbar_for_1_1_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_4_itm_1
          <= 1'b0;
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1 <= 1'b0;
      rva_in_reg_rw_sva_4 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_4
          <= 1'b0;
      GBCore_PushOutputs_switch_lp_asn_itm_3 <= 3'b000;
    end
    else if ( large_mem_write_arbxbar_xbar_for_1_for_and_cse ) begin
      large_mem_write_arbxbar_xbar_for_1_16_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[15];
      large_mem_write_arbxbar_xbar_for_1_15_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[14];
      large_mem_write_arbxbar_xbar_for_1_14_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[13];
      large_mem_write_arbxbar_xbar_for_1_13_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[12];
      large_mem_write_arbxbar_xbar_for_1_12_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[11];
      large_mem_write_arbxbar_xbar_for_1_11_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[10];
      large_mem_write_arbxbar_xbar_for_1_10_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[9];
      large_mem_write_arbxbar_xbar_for_1_9_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[8];
      large_mem_write_arbxbar_xbar_for_1_8_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[7];
      large_mem_write_arbxbar_xbar_for_1_7_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[6];
      large_mem_write_arbxbar_xbar_for_1_6_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[5];
      large_mem_write_arbxbar_xbar_for_1_5_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[4];
      large_mem_write_arbxbar_xbar_for_1_4_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[3];
      large_mem_write_arbxbar_xbar_for_1_3_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[2];
      large_mem_write_arbxbar_xbar_for_1_2_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_5_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[1];
      large_mem_write_arbxbar_xbar_for_1_1_for_large_mem_write_arbxbar_xbar_for_1_for_slc_large_mem_write_arbxbar_xbar_requests_transpose_1_0_4_itm_1
          <= large_mem_write_arbxbar_xbar_for_lshift_tmp[0];
      crossbar_spec_GB_Large_WordType_16U_16U_for_land_1_lpi_1_dfm_1 <= ~(crossbar_spec_GB_Large_WordType_16U_16U_for_mux_tmp
          | (~ large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_and_tmp));
      rva_in_reg_rw_sva_4 <= rva_in_reg_rw_sva_3;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_4
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
      GBCore_PushOutputs_switch_lp_asn_itm_3 <= GBCore_PushOutputs_switch_lp_asn_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_req_reg_is_write_sva_2 <= 1'b0;
      GBCore_SetLargeBuffer_1U_base_addr_acc_3_1 <= 16'b0000000000000000;
    end
    else if ( large_req_reg_is_write_and_cse ) begin
      large_req_reg_is_write_sva_2 <= large_req_reg_is_write_sva_1;
      GBCore_SetLargeBuffer_1U_base_addr_acc_3_1 <= GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_z;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_55 ) begin
      GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_15_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_32_enex5 ) begin
      large_write_data_data_0_15_lpi_1_dfm_4_2_16 <= large_write_data_data_0_15_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_14_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_33_enex5 ) begin
      large_write_data_data_0_14_lpi_1_dfm_4_2_16 <= large_write_data_data_0_14_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_13_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_34_enex5 ) begin
      large_write_data_data_0_13_lpi_1_dfm_4_2_16 <= large_write_data_data_0_13_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_12_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_35_enex5 ) begin
      large_write_data_data_0_12_lpi_1_dfm_4_2_16 <= large_write_data_data_0_12_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_11_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_36_enex5 ) begin
      large_write_data_data_0_11_lpi_1_dfm_4_2_16 <= large_write_data_data_0_11_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_10_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_37_enex5 ) begin
      large_write_data_data_0_10_lpi_1_dfm_4_2_16 <= large_write_data_data_0_10_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_9_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_38_enex5 ) begin
      large_write_data_data_0_9_lpi_1_dfm_4_2_16 <= large_write_data_data_0_9_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_8_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_39_enex5 ) begin
      large_write_data_data_0_8_lpi_1_dfm_4_2_16 <= large_write_data_data_0_8_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_7_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_40_enex5 ) begin
      large_write_data_data_0_7_lpi_1_dfm_4_2_16 <= large_write_data_data_0_7_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_6_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_41_enex5 ) begin
      large_write_data_data_0_6_lpi_1_dfm_4_2_16 <= large_write_data_data_0_6_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_5_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_42_enex5 ) begin
      large_write_data_data_0_5_lpi_1_dfm_4_2_16 <= large_write_data_data_0_5_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_4_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_43_enex5 ) begin
      large_write_data_data_0_4_lpi_1_dfm_4_2_16 <= large_write_data_data_0_4_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_3_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_44_enex5 ) begin
      large_write_data_data_0_3_lpi_1_dfm_4_2_16 <= large_write_data_data_0_3_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_2_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_45_enex5 ) begin
      large_write_data_data_0_2_lpi_1_dfm_4_2_16 <= large_write_data_data_0_2_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_1_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_46_enex5 ) begin
      large_write_data_data_0_1_lpi_1_dfm_4_2_16 <= large_write_data_data_0_1_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_write_data_data_0_0_lpi_1_dfm_4_2_16 <= 8'b00000000;
    end
    else if ( large_write_data_data_and_47_enex5 ) begin
      large_write_data_data_0_0_lpi_1_dfm_4_2_16 <= large_write_data_data_0_0_lpi_1_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_mux_11_itm_2 <= 1'b0;
      large_read_req_valid_0_lpi_1_dfm_3_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= 1'b0;
      GBCore_PushOutputs_switch_lp_asn_itm_2 <= 3'b000;
      rva_in_reg_rw_sva_3 <= 1'b0;
      GBCore_PushOutputs_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( large_write_data_data_and_cse ) begin
      while_mux_11_itm_2 <= while_mux_11_itm_1;
      large_read_req_valid_0_lpi_1_dfm_3_2 <= large_read_req_valid_0_lpi_1_dfm_3_1;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
      GBCore_PushOutputs_switch_lp_asn_itm_2 <= GBCore_PushOutputs_switch_lp_asn_itm_1;
      rva_in_reg_rw_sva_3 <= rva_in_reg_rw_sva_st_2;
      GBCore_PushOutputs_switch_lp_equal_tmp_2 <= GBCore_PushOutputs_switch_lp_equal_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_while_if_and_3_itm_3 <= 16'b0000000000000000;
    end
    else if ( while_if_and_25_enex5 ) begin
      while_if_while_if_and_3_itm_3 <= while_if_while_if_and_3_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_while_if_and_1_itm_3 <= 16'b0000000000000000;
    end
    else if ( while_if_and_26_enex5 ) begin
      while_if_while_if_and_1_itm_3 <= while_if_while_if_and_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_req_reg_vector_index_sva_1_1 <= 8'b00000000;
      large_req_reg_timestep_index_sva_1 <= 16'b0000000000000000;
      large_req_reg_is_write_sva_1 <= 1'b0;
    end
    else if ( large_req_reg_vector_index_and_cse ) begin
      large_req_reg_vector_index_sva_1_1 <= nmp_large_req_PopNB_mioi_data_vector_index_rsc_z_mxwt;
      large_req_reg_timestep_index_sva_1 <= nmp_large_req_PopNB_mioi_data_timestep_index_rsc_z_mxwt;
      large_req_reg_is_write_sva_1 <= nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_1
          <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_59 ) begin
      GBCore_PollNMPPort_Connections_InBlocking_spec_GB_Large_DataReq_Connections_SYN_PORT_PopNB_return_sva_st_1
          <= nmp_large_req_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= 1'b0;
      while_mux_11_itm_1 <= 1'b0;
      large_write_data_data_0_15_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_14_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_13_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_12_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_11_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_10_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_9_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_8_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_7_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_6_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_5_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_4_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_3_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_2_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_1_lpi_1_dfm_4_1 <= 8'b00000000;
      large_write_data_data_0_0_lpi_1_dfm_4_1 <= 8'b00000000;
      large_read_req_valid_0_lpi_1_dfm_3_1 <= 1'b0;
      GBCore_PushOutputs_switch_lp_asn_itm_1 <= 3'b000;
      rva_in_reg_rw_sva_st_2 <= 1'b0;
      GBCore_PushOutputs_switch_lp_equal_tmp_1 <= 1'b0;
    end
    else if ( while_if_and_3_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1;
      while_mux_11_itm_1 <= MUX_s_1_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_20_nl,
          while_if_while_if_and_5_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_15_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_21_nl,
          while_if_while_if_and_20_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_14_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_22_nl,
          while_if_while_if_and_19_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_13_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_23_nl,
          while_if_while_if_and_18_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_12_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_24_nl,
          while_if_while_if_and_17_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_11_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_25_nl,
          while_if_while_if_and_16_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_10_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_26_nl,
          while_if_while_if_and_15_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_9_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_27_nl,
          while_if_while_if_and_14_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_8_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_28_nl,
          while_if_while_if_and_13_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_7_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_29_nl,
          while_if_while_if_and_12_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_6_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_30_nl,
          while_if_while_if_and_11_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_5_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_31_nl,
          while_if_while_if_and_10_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_4_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_32_nl,
          while_if_while_if_and_9_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_3_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_33_nl,
          while_if_while_if_and_8_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_2_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_34_nl,
          while_if_while_if_and_7_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_1_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_35_nl,
          while_if_while_if_and_6_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_write_data_data_0_0_lpi_1_dfm_4_1 <= MUX_v_8_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_and_36_nl,
          while_if_while_if_and_5_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      large_read_req_valid_0_lpi_1_dfm_3_1 <= MUX_s_1_2_2(GBCore_PollNMPPort_GBCore_PollNMPPort_nor_1_nl,
          while_if_while_if_and_6_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1);
      GBCore_PushOutputs_switch_lp_asn_itm_1 <= GBCore_PushOutputs_switch_lp_asn_itm_1_mx0;
      rva_in_reg_rw_sva_st_2 <= rva_in_reg_rw_sva_1;
      GBCore_PushOutputs_switch_lp_equal_tmp_1 <= (GBCore_PushOutputs_switch_lp_asn_itm_1_mx0==3'b101);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1
          <= 1'b0;
      rva_in_reg_rw_sva_1 <= 1'b0;
    end
    else if ( while_if_and_4_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_1
          <= rva_in_large_PopNB_mioi_return_rsc_z_mxwt;
      rva_in_reg_rw_sva_1 <= rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104_lpi_1
          <= 8'b00000000;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112_lpi_1
          <= 8'b00000000;
      large_port_read_out_data_0_0_sva <= 8'b00000000;
    end
    else if ( and_286_cse ) begin
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_7_0_lpi_1_mx0;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_15_8_lp000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_23_16_l000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000002;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_39_32_l000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000002;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000002;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000002;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_l000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000002;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000002;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000002;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000002;
      crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112_lpi_1
          <= crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000002;
      large_port_read_out_data_0_0_sva <= large_port_read_out_data_0_0_sva_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_4 <= 1'b0;
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= 1'b0;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_15_cse ) begin
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_4 <= GBCore_DecodeAxiRead_switch_lp_nor_13_itm_3;
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_31_16_ftd
          <= 8'b00000000;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_29_enex5 ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_31_16_ftd
          <= reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_31_16_ftd_1
          <= 8'b00000000;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_30_enex5 ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_31_16_ftd_1
          <= reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_7_0
          <= 8'b00000000;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_31_enex5 ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_4_7_0
          <= GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_3_7_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_mem_write_arbxbar_xbar_for_empty_sva_1 <= 16'b0000000000000000;
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1 <= 4'b0000;
    end
    else if ( large_mem_write_arbxbar_xbar_for_empty_and_cse ) begin
      large_mem_write_arbxbar_xbar_for_empty_sva_1 <= large_mem_write_arbxbar_xbar_for_lshift_tmp;
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1 <= MUX_v_4_2_2(4'b0000,
          large_read_addrs_0_lpi_1_dfm_4_mx1_3_0, large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_large_mem_run_1_if_for_and_tmp);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_55_48_sva_dfm_1_4 <= 8'b00000000;
      rva_out_reg_data_1_63_56_sva_dfm_1_4 <= 8'b00000000;
      rva_out_reg_data_1_87_80_sva_dfm_1_4 <= 8'b00000000;
      rva_out_reg_data_1_95_88_sva_dfm_1_4 <= 8'b00000000;
      rva_out_reg_data_1_119_112_sva_dfm_1_4 <= 8'b00000000;
      rva_out_reg_data_1_127_120_sva_dfm_1_4 <= 8'b00000000;
      rva_out_reg_data_1_39_32_sva_dfm_1_4 <= 8'b00000000;
      rva_out_reg_data_1_71_64_sva_dfm_1_4 <= 8'b00000000;
      rva_out_reg_data_1_103_96_sva_dfm_1_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_1_cse ) begin
      rva_out_reg_data_1_55_48_sva_dfm_1_4 <= MUX_v_8_2_2(rva_out_reg_data_1_55_48_sva_dfm_1_3,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_l000001,
          and_dcpl_204);
      rva_out_reg_data_1_63_56_sva_dfm_1_4 <= MUX_v_8_2_2(rva_out_reg_data_1_63_56_sva_dfm_1_3,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_55_48_l000001,
          and_dcpl_204);
      rva_out_reg_data_1_87_80_sva_dfm_1_4 <= MUX_v_8_2_2(rva_out_reg_data_1_87_80_sva_dfm_1_3,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_l000001,
          and_dcpl_204);
      rva_out_reg_data_1_95_88_sva_dfm_1_4 <= MUX_v_8_2_2(rva_out_reg_data_1_95_88_sva_dfm_1_3,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_l000001,
          and_dcpl_204);
      rva_out_reg_data_1_119_112_sva_dfm_1_4 <= MUX_v_8_2_2(rva_out_reg_data_1_119_112_sva_dfm_1_3,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001,
          and_dcpl_204);
      rva_out_reg_data_1_127_120_sva_dfm_1_4 <= MUX_v_8_2_2(rva_out_reg_data_1_127_120_sva_dfm_1_3,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112000001,
          and_dcpl_204);
      rva_out_reg_data_1_39_32_sva_dfm_1_4 <= MUX_v_8_2_2(rva_out_reg_data_1_39_32_sva_dfm_1_3,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_31_24_l000001,
          and_dcpl_204);
      rva_out_reg_data_1_71_64_sva_dfm_1_4 <= MUX_v_8_2_2(rva_out_reg_data_1_71_64_sva_dfm_1_3,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_l000001,
          and_dcpl_204);
      rva_out_reg_data_1_103_96_sva_dfm_1_4 <= MUX_v_8_2_2(rva_out_reg_data_1_103_96_sva_dfm_1_3,
          crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_l000001,
          and_dcpl_204);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      num_vector_large_1_sva <= 8'b00000001;
      num_vector_large_2_sva <= 8'b00000001;
      num_vector_large_3_sva <= 8'b00000001;
    end
    else if ( and_334_cse ) begin
      num_vector_large_1_sva <= num_vector_large_1_sva_mx1;
      num_vector_large_2_sva <= num_vector_large_2_sva_mx1;
      num_vector_large_3_sva <= num_vector_large_3_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_4 <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_63 ) begin
      rva_in_reg_rw_sva_st_4 <= rva_in_reg_rw_sva_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_while_if_and_3_itm_2 <= 16'b0000000000000000;
    end
    else if ( while_if_and_27_enex5 ) begin
      while_if_while_if_and_3_itm_2 <= base_large_2_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_while_if_and_1_itm_2 <= 16'b0000000000000000;
    end
    else if ( while_if_and_28_enex5 ) begin
      while_if_while_if_and_1_itm_2 <= base_large_1_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      base_large_1_sva <= 16'b0000000000000000;
      base_large_2_sva <= 16'b0000000000000000;
    end
    else if ( base_large_and_cse ) begin
      base_large_1_sva <= MUX_v_16_2_2(base_large_1_sva_dfm_3_1, while_if_while_if_and_1_nl,
          and_cse);
      base_large_2_sva <= MUX_v_16_2_2(base_large_2_sva_dfm_3_1, while_if_while_if_and_3_nl,
          and_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      num_vector_large_3_sva_dfm_3_1 <= 8'b00000000;
      num_vector_large_2_sva_dfm_3_1 <= 8'b00000000;
      num_vector_large_1_sva_dfm_3_1 <= 8'b00000000;
      num_vector_large_0_sva_dfm_3_1 <= 8'b00000000;
      base_large_3_sva_dfm_3_1_15_8 <= 8'b00000000;
      base_large_3_sva_dfm_3_1_7_0 <= 8'b00000000;
      base_large_2_sva_dfm_3_1 <= 16'b0000000000000000;
      base_large_1_sva_dfm_3_1 <= 16'b0000000000000000;
      base_large_0_sva_dfm_3_1 <= 16'b0000000000000000;
    end
    else if ( and_363_cse ) begin
      num_vector_large_3_sva_dfm_3_1 <= MUX_v_8_2_2((rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[103:96]),
          num_vector_large_3_sva_mx1, or_dcpl_71);
      num_vector_large_2_sva_dfm_3_1 <= MUX_v_8_2_2((rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[71:64]),
          num_vector_large_2_sva_mx1, or_dcpl_71);
      num_vector_large_1_sva_dfm_3_1 <= MUX_v_8_2_2((rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[39:32]),
          num_vector_large_1_sva_mx1, or_dcpl_71);
      num_vector_large_0_sva_dfm_3_1 <= MUX_v_8_2_2((rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[7:0]),
          num_vector_large_0_sva_mx0, or_dcpl_71);
      base_large_3_sva_dfm_3_1_15_8 <= MUX_v_8_2_2((rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[127:120]),
          base_large_3_sva_mx2_15_8, or_dcpl_71);
      base_large_3_sva_dfm_3_1_7_0 <= MUX_v_8_2_2((rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[119:112]),
          base_large_3_sva_mx2_7_0, or_dcpl_71);
      base_large_2_sva_dfm_3_1 <= MUX_v_16_2_2((rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[95:80]),
          base_large_2_sva_mx1, or_dcpl_71);
      base_large_1_sva_dfm_3_1 <= MUX_v_16_2_2((rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[63:48]),
          base_large_1_sva_mx1, or_dcpl_71);
      base_large_0_sva_dfm_3_1 <= MUX_v_16_2_2((rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[31:16]),
          base_large_0_sva_mx0, or_dcpl_71);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_while_if_and_20_itm_1 <= 8'b00000000;
      while_if_while_if_and_19_itm_1 <= 8'b00000000;
      while_if_while_if_and_18_itm_1 <= 8'b00000000;
      while_if_while_if_and_17_itm_1 <= 8'b00000000;
      while_if_while_if_and_16_itm_1 <= 8'b00000000;
      while_if_while_if_and_15_itm_1 <= 8'b00000000;
      while_if_while_if_and_14_itm_1 <= 8'b00000000;
      while_if_while_if_and_13_itm_1 <= 8'b00000000;
      while_if_while_if_and_12_itm_1 <= 8'b00000000;
      while_if_while_if_and_11_itm_1 <= 8'b00000000;
      while_if_while_if_and_10_itm_1 <= 8'b00000000;
      while_if_while_if_and_9_itm_1 <= 8'b00000000;
      while_if_while_if_and_8_itm_1 <= 8'b00000000;
      while_if_while_if_and_7_itm_1 <= 8'b00000000;
      while_if_while_if_and_6_itm_1 <= 8'b00000000;
      while_if_while_if_and_5_itm_1 <= 8'b00000000;
      while_if_while_if_and_itm_1 <= 3'b000;
    end
    else if ( while_if_and_8_cse ) begin
      while_if_while_if_and_20_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[127:120])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_19_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[119:112])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_18_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[111:104])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_17_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[103:96])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_16_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[95:88])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_15_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[87:80])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_14_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[79:72])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_13_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[71:64])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_12_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[63:56])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_11_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[55:48])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_10_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[47:40])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_9_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[39:32])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_8_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[31:24])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_7_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[23:16])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_6_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[15:8])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_5_itm_1 <= (rva_in_large_PopNB_mioi_data_data_rsc_z_mxwt[7:0])
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0})
          & ({{7{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt});
      while_if_while_if_and_itm_1 <= ~(GBCore_DecodeAxiRead_switch_lp_mux1h_20_nl
          | ({{2{GBCore_DecodeAxiRead_switch_lp_nor_tmp_1}}, GBCore_DecodeAxiRead_switch_lp_nor_tmp_1})
          | ({{2{rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_3 <= 1'b0;
    end
    else if ( while_if_and_cse ) begin
      rva_in_reg_rw_sva_st_3 <= rva_in_reg_rw_sva_st_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_3 <= 1'b0;
    end
    else if ( GBCoreRun_wen & and_dcpl_58 & (~ rva_in_reg_rw_sva_st_2) ) begin
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_3 <= GBCore_DecodeAxiRead_switch_lp_nor_13_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_3_7_0
          <= 8'b00000000;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_20_enex5 ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_3_7_0
          <= GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_7_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_103_96_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_54_enex5 ) begin
      rva_out_reg_data_1_103_96_sva_dfm_1_3 <= rva_out_reg_data_1_103_96_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_71_64_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_55_enex5 ) begin
      rva_out_reg_data_1_71_64_sva_dfm_1_3 <= rva_out_reg_data_1_71_64_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_39_32_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_56_enex5 ) begin
      rva_out_reg_data_1_39_32_sva_dfm_1_3 <= rva_out_reg_data_1_39_32_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_127_120_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_57_enex5 ) begin
      rva_out_reg_data_1_127_120_sva_dfm_1_3 <= rva_out_reg_data_1_127_120_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_119_112_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_58_enex5 ) begin
      rva_out_reg_data_1_119_112_sva_dfm_1_3 <= rva_out_reg_data_1_119_112_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_95_88_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_59_enex5 ) begin
      rva_out_reg_data_1_95_88_sva_dfm_1_3 <= rva_out_reg_data_1_95_88_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_87_80_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_60_enex5 ) begin
      rva_out_reg_data_1_87_80_sva_dfm_1_3 <= rva_out_reg_data_1_87_80_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_63_56_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_61_enex5 ) begin
      rva_out_reg_data_1_63_56_sva_dfm_1_3 <= rva_out_reg_data_1_63_56_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_55_48_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_62_enex5 ) begin
      rva_out_reg_data_1_55_48_sva_dfm_1_3 <= rva_out_reg_data_1_55_48_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( GBCoreRun_wen & (~(nand_17_cse | (~ rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt)))
        ) begin
      GBCore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_3 <= 1'b0;
    end
    else if ( GBCoreRun_wen & (~(nand_17_cse | rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt))
        ) begin
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_3 <= GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_2 <= 1'b0;
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_21_cse ) begin
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_2 <= GBCore_DecodeAxiRead_switch_lp_nor_13_itm_1;
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_7_0
          <= 8'b00000000;
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_24
          <= 8'b00000000;
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_23_16
          <= 8'b00000000;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_23_cse ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_7_0
          <= MUX1HOT_v_8_4_2(GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_7_0,
          num_vector_large_1_sva, num_vector_large_2_sva, num_vector_large_3_sva,
          {GBCore_DecodeAxiRead_switch_lp_or_4_cse , GBCore_DecodeAxiRead_switch_lp_and_6_cse
          , GBCore_DecodeAxiRead_switch_lp_and_7_cse , GBCore_DecodeAxiRead_switch_lp_and_8_cse});
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_24
          <= MUX1HOT_v_8_4_2((GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_31_16[15:8]),
          (base_large_1_sva[15:8]), (base_large_2_sva[15:8]), base_large_3_sva_15_8,
          {GBCore_DecodeAxiRead_switch_lp_or_4_cse , GBCore_DecodeAxiRead_switch_lp_and_6_cse
          , GBCore_DecodeAxiRead_switch_lp_and_7_cse , GBCore_DecodeAxiRead_switch_lp_and_8_cse});
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_23_16
          <= MUX1HOT_v_8_4_2((GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_31_16[7:0]),
          (base_large_1_sva[7:0]), (base_large_2_sva[7:0]), base_large_3_sva_7_0,
          {GBCore_DecodeAxiRead_switch_lp_or_4_cse , GBCore_DecodeAxiRead_switch_lp_and_6_cse
          , GBCore_DecodeAxiRead_switch_lp_and_7_cse , GBCore_DecodeAxiRead_switch_lp_and_8_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_103_96_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_63_enex5 ) begin
      rva_out_reg_data_1_103_96_sva_dfm_1_2 <= base_large_3_sva_7_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_71_64_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_64_enex5 ) begin
      rva_out_reg_data_1_71_64_sva_dfm_1_2 <= rva_out_reg_data_1_71_64_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_39_32_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_65_enex5 ) begin
      rva_out_reg_data_1_39_32_sva_dfm_1_2 <= rva_out_reg_data_1_39_32_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_127_120_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_66_enex5 ) begin
      rva_out_reg_data_1_127_120_sva_dfm_1_2 <= rva_out_reg_data_1_127_120_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_119_112_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_67_enex5 ) begin
      rva_out_reg_data_1_119_112_sva_dfm_1_2 <= rva_out_reg_data_1_119_112_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_95_88_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_68_enex5 ) begin
      rva_out_reg_data_1_95_88_sva_dfm_1_2 <= rva_out_reg_data_1_95_88_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_87_80_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_69_enex5 ) begin
      rva_out_reg_data_1_87_80_sva_dfm_1_2 <= rva_out_reg_data_1_87_80_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_63_56_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_70_enex5 ) begin
      rva_out_reg_data_1_63_56_sva_dfm_1_2 <= rva_out_reg_data_1_63_56_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_1_55_48_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_71_enex5 ) begin
      rva_out_reg_data_1_55_48_sva_dfm_1_2 <= rva_out_reg_data_1_55_48_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_1 <= 1'b0;
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= 1'b0;
      rva_out_reg_data_1_71_64_sva_dfm_1_1 <= 8'b00000000;
      rva_out_reg_data_1_39_32_sva_dfm_1_1 <= 8'b00000000;
      rva_out_reg_data_1_127_120_sva_dfm_1_1 <= 8'b00000000;
      rva_out_reg_data_1_119_112_sva_dfm_1_1 <= 8'b00000000;
      rva_out_reg_data_1_95_88_sva_dfm_1_1 <= 8'b00000000;
      rva_out_reg_data_1_87_80_sva_dfm_1_1 <= 8'b00000000;
      rva_out_reg_data_1_63_56_sva_dfm_1_1 <= 8'b00000000;
      rva_out_reg_data_1_55_48_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_25_cse ) begin
      GBCore_DecodeAxiRead_switch_lp_nor_13_itm_1 <= ~(GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          | GBCore_DecodeAxiRead_switch_lp_nor_tmp_1);
      GBCore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= GBCore_DecodeAxiRead_switch_lp_equal_tmp_4;
      rva_out_reg_data_1_71_64_sva_dfm_1_1 <= num_vector_large_2_sva_mx1 & (signext_8_1(~
          GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse))
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_4}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_4});
      rva_out_reg_data_1_39_32_sva_dfm_1_1 <= num_vector_large_1_sva_mx1 & (signext_8_1(~
          GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse))
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_4}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_4});
      rva_out_reg_data_1_127_120_sva_dfm_1_1 <= base_large_3_sva_mx2_15_8 & (signext_8_1(~
          GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse))
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_4}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_4});
      rva_out_reg_data_1_119_112_sva_dfm_1_1 <= base_large_3_sva_mx2_7_0 & (signext_8_1(~
          GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse))
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_4}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_4});
      rva_out_reg_data_1_95_88_sva_dfm_1_1 <= (base_large_2_sva_mx1[15:8]) & (signext_8_1(~
          GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse))
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_4}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_4});
      rva_out_reg_data_1_87_80_sva_dfm_1_1 <= (base_large_2_sva_mx1[7:0]) & (signext_8_1(~
          GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse))
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_4}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_4});
      rva_out_reg_data_1_63_56_sva_dfm_1_1 <= (base_large_1_sva_mx1[15:8]) & (signext_8_1(~
          GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse))
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_4}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_4});
      rva_out_reg_data_1_55_48_sva_dfm_1_1 <= (base_large_1_sva_mx1[7:0]) & (signext_8_1(~
          GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse))
          & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_4}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_4});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_31_16
          <= 16'b0000000000000000;
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_7_0
          <= 8'b00000001;
    end
    else if ( and_549_cse ) begin
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_31_16
          <= MUX_v_16_2_2(GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_21_nl,
          base_large_0_sva_dfm_3_1, and_dcpl_206);
      GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_1_7_0
          <= MUX_v_8_2_2(GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_20_nl,
          num_vector_large_0_sva_dfm_3_1, and_dcpl_206);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_0 <= 8'b00000000;
    end
    else if ( GBCore_SetLargeBuffer_1U_base_addr_and_2_enex5 ) begin
      reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_0 <= GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_24;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_1 <= 8'b00000000;
    end
    else if ( GBCore_SetLargeBuffer_1U_base_addr_and_3_enex5 ) begin
      reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_cse_rsp_1 <= GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_23_16;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      base_large_3_sva_15_8 <= 8'b00000000;
    end
    else if ( base_large_and_8_enex5 ) begin
      base_large_3_sva_15_8 <= base_large_3_sva_dfm_3_1_15_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      base_large_3_sva_7_0 <= 8'b00000000;
    end
    else if ( base_large_and_3_ssc ) begin
      base_large_3_sva_7_0 <= MUX_v_8_2_2(base_large_3_sva_dfm_3_1_7_0, GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_7_nl,
          and_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_127_120_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_45_enex5 ) begin
      reg_rva_out_reg_data_1_127_120_sva_dfm_1_4_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_119_112_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_46_enex5 ) begin
      reg_rva_out_reg_data_1_119_112_sva_dfm_1_4_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_103_96_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_47_enex5 ) begin
      reg_rva_out_reg_data_1_103_96_sva_dfm_1_4_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_95_88_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_48_enex5 ) begin
      reg_rva_out_reg_data_1_95_88_sva_dfm_1_4_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_39_32_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_49_enex5 ) begin
      reg_rva_out_reg_data_1_39_32_sva_dfm_1_4_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_87_80_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_50_enex5 ) begin
      reg_rva_out_reg_data_1_87_80_sva_dfm_1_4_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_55_48_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_51_enex5 ) begin
      reg_rva_out_reg_data_1_55_48_sva_dfm_1_4_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_71_64_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_52_enex5 ) begin
      reg_rva_out_reg_data_1_71_64_sva_dfm_1_4_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_63_56_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_53_enex5 ) begin
      reg_rva_out_reg_data_1_63_56_sva_dfm_1_4_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_15_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_32_enex5 ) begin
      reg_large_write_data_data_0_15_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_14_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_33_enex5 ) begin
      reg_large_write_data_data_0_14_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_13_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_34_enex5 ) begin
      reg_large_write_data_data_0_13_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_12_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_35_enex5 ) begin
      reg_large_write_data_data_0_12_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_11_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_36_enex5 ) begin
      reg_large_write_data_data_0_11_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_10_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_37_enex5 ) begin
      reg_large_write_data_data_0_10_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_9_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_38_enex5 ) begin
      reg_large_write_data_data_0_9_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_8_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_39_enex5 ) begin
      reg_large_write_data_data_0_8_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_7_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_40_enex5 ) begin
      reg_large_write_data_data_0_7_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_6_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_41_enex5 ) begin
      reg_large_write_data_data_0_6_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_5_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_42_enex5 ) begin
      reg_large_write_data_data_0_5_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_4_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_43_enex5 ) begin
      reg_large_write_data_data_0_4_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_3_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_44_enex5 ) begin
      reg_large_write_data_data_0_3_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_2_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_45_enex5 ) begin
      reg_large_write_data_data_0_2_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_1_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_46_enex5 ) begin
      reg_large_write_data_data_0_1_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_large_write_data_data_0_0_lpi_1_dfm_4_1_enexo <= 1'b1;
    end
    else if ( while_if_and_3_cse | large_write_data_data_and_47_enex5 ) begin
      reg_large_write_data_data_0_0_lpi_1_dfm_4_1_enexo <= while_if_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_if_while_if_and_3_itm_2_enexo <= 1'b1;
    end
    else if ( while_if_and_27_enex5 | while_if_and_25_enex5 ) begin
      reg_while_if_while_if_and_3_itm_2_enexo <= while_if_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_if_while_if_and_1_itm_2_enexo <= 1'b1;
    end
    else if ( while_if_and_28_enex5 | while_if_and_26_enex5 ) begin
      reg_while_if_while_if_and_1_itm_2_enexo <= while_if_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_enexo <= 1'b1;
    end
    else if ( GBCore_SetLargeBuffer_1U_base_addr_and_2_enex5 | GBCore_DecodeAxiRead_switch_lp_and_29_enex5
        ) begin
      reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_enexo <= GBCore_SetLargeBuffer_1U_base_addr_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_1_enexo <= 1'b1;
    end
    else if ( GBCore_SetLargeBuffer_1U_base_addr_and_3_enex5 | GBCore_DecodeAxiRead_switch_lp_and_30_enex5
        ) begin
      reg_GBCore_SetLargeBuffer_1U_base_addr_mux_itm_2_1_enexo <= GBCore_SetLargeBuffer_1U_base_addr_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_3_7_0_enexo
          <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_20_enex5 | GBCore_DecodeAxiRead_switch_lp_and_31_enex5
        ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_3_7_0_enexo
          <= GBCore_DecodeAxiRead_switch_lp_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_base_large_2_enexo <= 1'b1;
    end
    else if ( base_large_and_cse | while_if_and_27_enex5 ) begin
      reg_base_large_2_enexo <= base_large_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_base_large_1_enexo <= 1'b1;
    end
    else if ( base_large_and_cse | while_if_and_28_enex5 ) begin
      reg_base_large_1_enexo <= base_large_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_7_0_enexo
          <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_23_cse | GBCore_DecodeAxiRead_switch_lp_and_20_enex5
        ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_7_0_enexo
          <= GBCore_DecodeAxiRead_switch_lp_and_23_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_103_96_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_63_enex5 | rva_out_reg_data_and_54_enex5 ) begin
      reg_rva_out_reg_data_1_103_96_sva_dfm_1_2_enexo <= rva_out_reg_data_and_63_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_71_64_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_64_enex5 | rva_out_reg_data_and_55_enex5 ) begin
      reg_rva_out_reg_data_1_71_64_sva_dfm_1_2_enexo <= rva_out_reg_data_and_64_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_39_32_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_65_enex5 | rva_out_reg_data_and_56_enex5 ) begin
      reg_rva_out_reg_data_1_39_32_sva_dfm_1_2_enexo <= rva_out_reg_data_and_65_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_127_120_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_66_enex5 | rva_out_reg_data_and_57_enex5 ) begin
      reg_rva_out_reg_data_1_127_120_sva_dfm_1_2_enexo <= rva_out_reg_data_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_119_112_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_67_enex5 | rva_out_reg_data_and_58_enex5 ) begin
      reg_rva_out_reg_data_1_119_112_sva_dfm_1_2_enexo <= rva_out_reg_data_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_95_88_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_68_enex5 | rva_out_reg_data_and_59_enex5 ) begin
      reg_rva_out_reg_data_1_95_88_sva_dfm_1_2_enexo <= rva_out_reg_data_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_87_80_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_69_enex5 | rva_out_reg_data_and_60_enex5 ) begin
      reg_rva_out_reg_data_1_87_80_sva_dfm_1_2_enexo <= rva_out_reg_data_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_63_56_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_70_enex5 | rva_out_reg_data_and_61_enex5 ) begin
      reg_rva_out_reg_data_1_63_56_sva_dfm_1_2_enexo <= rva_out_reg_data_and_70_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_55_48_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_71_enex5 | rva_out_reg_data_and_62_enex5 ) begin
      reg_rva_out_reg_data_1_55_48_sva_dfm_1_2_enexo <= rva_out_reg_data_and_71_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_base_large_3_1_enexo <= 1'b1;
    end
    else if ( base_large_and_3_ssc | rva_out_reg_data_and_63_enex5 ) begin
      reg_base_large_3_1_enexo <= base_large_and_3_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_71_64_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_25_cse | rva_out_reg_data_and_64_enex5
        ) begin
      reg_rva_out_reg_data_1_71_64_sva_dfm_1_1_enexo <= GBCore_DecodeAxiRead_switch_lp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_39_32_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_25_cse | rva_out_reg_data_and_65_enex5
        ) begin
      reg_rva_out_reg_data_1_39_32_sva_dfm_1_1_enexo <= GBCore_DecodeAxiRead_switch_lp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_127_120_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_25_cse | rva_out_reg_data_and_66_enex5
        ) begin
      reg_rva_out_reg_data_1_127_120_sva_dfm_1_1_enexo <= GBCore_DecodeAxiRead_switch_lp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_119_112_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_25_cse | rva_out_reg_data_and_67_enex5
        ) begin
      reg_rva_out_reg_data_1_119_112_sva_dfm_1_1_enexo <= GBCore_DecodeAxiRead_switch_lp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_95_88_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_25_cse | rva_out_reg_data_and_68_enex5
        ) begin
      reg_rva_out_reg_data_1_95_88_sva_dfm_1_1_enexo <= GBCore_DecodeAxiRead_switch_lp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_87_80_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_25_cse | rva_out_reg_data_and_69_enex5
        ) begin
      reg_rva_out_reg_data_1_87_80_sva_dfm_1_1_enexo <= GBCore_DecodeAxiRead_switch_lp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_63_56_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_25_cse | rva_out_reg_data_and_70_enex5
        ) begin
      reg_rva_out_reg_data_1_63_56_sva_dfm_1_1_enexo <= GBCore_DecodeAxiRead_switch_lp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_1_55_48_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_25_cse | rva_out_reg_data_and_71_enex5
        ) begin
      reg_rva_out_reg_data_1_55_48_sva_dfm_1_1_enexo <= GBCore_DecodeAxiRead_switch_lp_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_16_enexo
          <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_23_cse | GBCore_SetLargeBuffer_1U_base_addr_and_2_enex5
        ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_16_enexo
          <= GBCore_DecodeAxiRead_switch_lp_and_23_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_16_1_enexo
          <= 1'b1;
    end
    else if ( GBCore_DecodeAxiRead_switch_lp_and_23_cse | GBCore_SetLargeBuffer_1U_base_addr_and_3_enex5
        ) begin
      reg_GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_10_itm_2_31_16_1_enexo
          <= GBCore_DecodeAxiRead_switch_lp_and_23_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_base_large_3_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( and_363_cse | base_large_and_8_enex5 ) begin
      reg_base_large_3_sva_dfm_3_1_enexo <= and_363_cse;
    end
  end
  assign or_85_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | rva_in_reg_rw_sva_st_2 | (~ while_stage_0_4);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_262_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_262_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_264_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_16_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_264_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_266_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_32_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_266_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_268_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_48_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_268_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_270_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_64_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_270_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_272_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_80_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_272_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_274_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_96_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_274_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_276_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_112_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_276_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_278_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_128_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_278_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_280_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_144_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_280_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_282_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_160_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_282_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_284_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_176_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_284_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_286_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_192_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_286_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_256_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_208_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_256_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_258_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_224_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_258_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_260_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_240_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[7:0]),
      large_mem_write_arbxbar_xbar_for_1_for_not_260_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_1_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_o000000
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_16_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_32_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_48_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_64_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_80_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_96_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_112_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_128_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_144_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_160_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_176_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_192_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_208_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_224_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_240_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_333_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_1_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_333_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_348_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_17_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_348_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_363_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_33_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_363_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_378_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_49_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_378_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_393_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_65_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_393_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_408_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_81_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_408_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_423_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_97_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_423_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_438_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_113_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_438_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_453_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_129_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_453_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_468_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_145_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_468_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_483_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_161_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_483_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_498_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_177_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_498_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_513_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_193_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_513_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_288_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_209_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_288_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_303_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_225_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_303_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_318_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_241_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[15:8]),
      large_mem_write_arbxbar_xbar_for_1_for_not_318_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000000
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_1_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_17_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_33_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_49_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_65_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_81_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_97_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_113_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_129_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_145_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_161_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_177_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_193_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_209_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_225_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_241_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_345_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_13_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_345_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_360_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_29_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_360_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_375_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_45_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_375_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_390_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_61_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_390_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_405_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_77_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_405_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_420_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_93_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_420_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_435_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_109_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_435_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_450_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_125_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_450_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_465_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_141_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_465_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_480_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_157_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_480_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_495_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_173_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_495_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_510_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_189_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_510_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_525_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_205_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_525_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_300_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_221_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_300_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_315_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_237_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_315_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_330_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_253_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[111:104]),
      large_mem_write_arbxbar_xbar_for_1_for_not_330_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000001
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_13_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_29_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_45_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_61_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_77_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_93_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_109_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_125_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_141_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_157_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_173_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_189_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_205_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_221_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_237_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_253_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_334_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_2_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_334_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_349_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_18_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_349_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_364_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_34_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_364_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_379_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_50_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_379_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_394_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_66_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_394_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_409_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_82_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_409_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_424_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_98_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_424_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_439_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_114_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_439_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_454_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_130_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_454_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_469_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_146_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_469_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_484_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_162_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_484_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_499_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_178_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_499_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_514_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_194_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_514_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_289_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_210_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_289_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_304_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_226_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_304_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_319_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_242_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[23:16]),
      large_mem_write_arbxbar_xbar_for_1_for_not_319_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000002
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_2_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_18_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_34_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_50_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_66_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_82_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_98_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_114_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_130_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_146_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_162_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_178_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_194_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_210_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_226_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_242_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_335_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_3_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_335_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_350_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_19_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_350_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_365_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_35_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_365_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_380_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_51_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_380_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_395_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_67_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_395_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_410_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_83_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_410_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_425_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_99_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_425_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_440_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_115_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_440_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_455_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_131_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_455_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_470_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_147_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_470_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_485_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_163_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_485_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_500_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_179_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_500_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_515_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_195_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_515_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_290_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_211_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_290_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_305_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_227_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_305_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_320_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_243_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[31:24]),
      large_mem_write_arbxbar_xbar_for_1_for_not_320_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000003
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_3_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_19_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_35_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_51_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_67_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_83_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_99_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_115_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_131_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_147_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_163_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_179_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_195_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_211_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_227_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_243_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_337_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_5_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_337_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_352_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_21_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_352_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_367_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_37_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_367_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_382_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_53_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_382_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_397_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_69_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_397_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_412_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_85_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_412_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_427_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_101_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_427_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_442_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_117_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_442_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_457_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_133_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_457_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_472_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_149_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_472_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_487_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_165_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_487_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_502_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_181_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_502_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_517_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_197_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_517_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_292_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_213_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_292_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_307_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_229_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_307_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_322_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_245_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[47:40]),
      large_mem_write_arbxbar_xbar_for_1_for_not_322_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000004
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_5_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_21_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_37_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_53_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_69_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_85_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_101_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_117_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_133_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_149_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_165_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_181_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_197_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_213_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_229_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_245_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_341_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[0]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_9_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_341_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_356_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[1]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_25_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_356_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_371_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_41_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_371_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_386_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_57_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_386_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_401_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_73_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_401_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_416_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_89_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_416_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_431_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_105_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_431_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_446_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_121_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_446_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_461_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[8]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_137_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_461_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_476_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[9]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_153_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_476_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_491_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[10]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_169_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_491_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_506_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[11]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_185_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_506_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_521_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[12]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_201_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_521_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_296_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[13]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_217_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_296_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_311_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[14]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_233_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_311_nl);
  assign large_mem_write_arbxbar_xbar_for_1_for_not_326_nl = ~ (large_mem_write_arbxbar_xbar_for_empty_sva_1[15]);
  assign large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_249_nl
      = MUX_v_8_2_2(8'b00000000, (large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d[79:72]),
      large_mem_write_arbxbar_xbar_for_1_for_not_326_nl);
  assign crossbar_spec_GB_Large_WordType_16U_16U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_large_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_data_in_tmp_000005
      = MUX_v_8_16_2(large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_9_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_25_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_41_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_57_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_73_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_89_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_105_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_121_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_137_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_153_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_169_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_185_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_201_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_217_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_233_nl,
      large_mem_banks_load_store_for_else_large_mem_banks_load_store_for_else_and_249_nl,
      crossbar_spec_GB_Large_WordType_16U_16U_source_tmp_1_lpi_1_dfm_1);
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_20_nl = nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt
      & nmp_large_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_if_while_if_and_5_nl = GBCore_DecodeAxiWrite_switch_lp_equal_tmp_2
      & rva_in_reg_rw_sva_1;
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_21_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[127:120])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_22_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[119:112])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_23_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[111:104])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_24_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[103:96])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_25_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[95:88])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_26_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[87:80])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_27_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[79:72])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_28_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[71:64])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_29_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[63:56])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_30_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[55:48])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_31_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[47:40])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_32_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[39:32])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_33_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[31:24])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_34_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[23:16])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_35_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[15:8])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_and_36_nl = (nmp_large_req_PopNB_mioi_data_write_data_data_rsc_z_mxwt[7:0])
      & ({{7{nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt})
      & ({{7{nmp_large_req_PopNB_mioi_return_rsc_z_mxwt}}, nmp_large_req_PopNB_mioi_return_rsc_z_mxwt});
  assign GBCore_PollNMPPort_GBCore_PollNMPPort_nor_1_nl = ~(nmp_large_req_PopNB_mioi_data_is_write_rsc_z_mxwt
      | (~ nmp_large_req_PopNB_mioi_return_rsc_z_mxwt));
  assign while_if_while_if_and_6_nl = GBCore_DecodeAxiRead_switch_lp_equal_tmp_3
      & (~ rva_in_reg_rw_sva_1);
  assign rva_in_reg_rw_not_42_nl = ~ rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign while_if_while_if_and_1_nl = MUX_v_16_2_2(16'b0000000000000000, large_write_addrs_lpi_1_dfm_6,
      rva_in_reg_rw_not_42_nl);
  assign while_if_while_if_and_3_nl = MUX_v_16_2_2(16'b0000000000000000, large_write_addrs_lpi_1_dfm_6,
      rva_in_large_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign GBCore_DecodeAxiRead_switch_lp_mux1h_20_nl = MUX1HOT_v_3_3_2(3'b100, 3'b011,
      3'b010, {GBCore_DecodeAxiRead_switch_lp_equal_tmp_5 , GBCore_DecodeAxiRead_switch_lp_equal_tmp_4
      , GBCore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0});
  assign GBCore_DecodeAxiRead_switch_lp_not_20_nl = ~ GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse;
  assign GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_21_nl
      = MUX_v_16_2_2(16'b0000000000000000, base_large_0_sva_mx0, GBCore_DecodeAxiRead_switch_lp_not_20_nl);
  assign GBCore_DecodeAxiRead_switch_lp_not_19_nl = ~ GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse;
  assign GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_20_nl
      = MUX_v_8_2_2(8'b00000000, num_vector_large_0_sva_mx0, GBCore_DecodeAxiRead_switch_lp_not_19_nl);
  assign GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_and_7_nl =
      num_vector_large_3_sva_mx1 & (signext_8_1(~ GBCore_DecodeAxiRead_switch_lp_GBCore_DecodeAxiRead_switch_lp_nand_cse))
      & ({{7{GBCore_DecodeAxiRead_switch_lp_equal_tmp_4}}, GBCore_DecodeAxiRead_switch_lp_equal_tmp_4});

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_16_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input  input_8;
    input  input_9;
    input  input_10;
    input  input_11;
    input  input_12;
    input  input_13;
    input  input_14;
    input  input_15;
    input [3:0] sel;
    reg  result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_s_1_16_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input  sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_16_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [3:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_8_16_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [15:0] signext_16_1;
    input  vector;
  begin
    signext_16_1= {{15{vector}}, vector};
  end
  endfunction


  function automatic [7:0] signext_8_1;
    input  vector;
  begin
    signext_8_1= {{7{vector}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP_NMPRun
// ------------------------------------------------------------------


module GBModule_NMP_NMPRun (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      start_vld, start_rdy, start_dat, done_vld, done_rdy, done_dat, large_req_vld,
      large_req_rdy, large_req_dat, large_rsp_vld, large_rsp_rdy, large_rsp_dat,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_a, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_z, NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_a,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_z, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_b,
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_a, NMP_ComputeRMSNormalize_for_1_mul_cmp_en,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_1_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_1_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_2_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_2_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_3_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_3_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_4_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_4_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_5_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_5_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_6_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_6_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_7_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_7_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_8_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_8_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_9_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_9_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_10_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_10_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_11_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_11_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_12_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_12_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_13_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_13_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_14_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_14_z, NMP_ComputeRMSNormalize_for_1_mul_cmp_15_a,
      NMP_ComputeRMSNormalize_for_1_mul_cmp_15_z, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_z, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_z,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_z, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_z,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_z, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_z,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_z, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_z,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_z, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_z,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_z, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_z,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_z, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_z,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_z, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_z,
      NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_pff, NMP_ComputeRMSNormalize_for_1_mul_cmp_b_pff,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_a_pff, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_a_pff,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_a_pff, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_a_pff,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_a_pff, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_a_pff,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_a_pff, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_a_pff,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_a_pff, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_a_pff,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_a_pff, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_a_pff,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_a_pff, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_a_pff,
      NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_a_pff, NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_a_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  input start_vld;
  output start_rdy;
  input start_dat;
  output done_vld;
  input done_rdy;
  output done_dat;
  output large_req_vld;
  input large_req_rdy;
  output [154:0] large_req_dat;
  input large_rsp_vld;
  output large_rsp_rdy;
  input [127:0] large_rsp_dat;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_a;
  output NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_z;
  output [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_a;
  input [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_b;
  output NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z;
  output [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_b;
  input [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_a;
  output NMP_ComputeRMSNormalize_for_1_mul_cmp_en;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_1_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_1_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_2_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_2_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_3_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_3_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_4_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_4_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_5_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_5_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_6_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_6_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_7_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_7_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_8_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_8_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_9_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_9_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_10_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_10_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_11_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_11_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_12_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_12_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_13_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_13_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_14_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_14_z;
  output [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_15_a;
  input [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_15_z;
  output NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_z;
  input [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_z;
  output [39:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_pff;
  output [39:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_b_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_a_pff;
  output [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_a_pff;


  // Interconnect Declarations
  wire NMPRun_wen;
  wire NMPRun_wten;
  wire [33:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire large_req_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire [127:0] large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt;
  wire large_rsp_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire done_Push_mioi_wen_comp;
  wire fsm_output;
  wire NMP_RunFSM_switch_lp_or_73_tmp;
  wire [39:0] operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_1_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_2_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_3_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_4_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_5_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_6_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_7_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_8_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_9_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_10_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_11_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_12_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_13_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_14_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_15_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_1_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_2_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_3_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_4_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_5_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_6_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_7_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_8_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_9_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_10_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_11_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_12_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_13_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_14_tmp;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_15_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp;
  wire [6:0] NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp;
  wire [7:0] nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp;
  wire NMP_ComputeSoftmaxMax_for_if_less_5_tmp;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_2;
  wire NMP_ComputeSoftmaxMax_for_if_less_12_tmp;
  wire nmp_config_ConfigRead_nor_2_tmp;
  wire and_dcpl;
  wire and_dcpl_3;
  wire and_dcpl_5;
  wire and_dcpl_6;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_10;
  wire or_dcpl_5;
  wire or_dcpl_12;
  wire or_dcpl_19;
  wire or_dcpl_26;
  wire or_dcpl_33;
  wire or_dcpl_40;
  wire or_dcpl_47;
  wire or_dcpl_54;
  wire or_dcpl_61;
  wire or_dcpl_68;
  wire or_dcpl_75;
  wire or_dcpl_82;
  wire or_dcpl_89;
  wire or_dcpl_96;
  wire or_dcpl_103;
  wire or_dcpl_110;
  wire and_dcpl_46;
  wire and_dcpl_47;
  wire or_dcpl_117;
  wire or_dcpl_124;
  wire or_dcpl_131;
  wire or_dcpl_138;
  wire or_dcpl_145;
  wire or_dcpl_152;
  wire or_dcpl_159;
  wire or_dcpl_166;
  wire or_dcpl_173;
  wire or_dcpl_180;
  wire or_dcpl_187;
  wire or_dcpl_194;
  wire or_dcpl_201;
  wire or_dcpl_208;
  wire or_dcpl_215;
  wire or_dcpl_222;
  wire and_dcpl_88;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_100;
  wire and_dcpl_101;
  wire and_dcpl_105;
  wire and_dcpl_108;
  wire and_dcpl_122;
  wire and_dcpl_124;
  wire and_dcpl_125;
  wire and_dcpl_129;
  wire and_dcpl_130;
  wire and_dcpl_134;
  wire and_dcpl_136;
  wire and_dcpl_137;
  wire and_dcpl_139;
  wire and_dcpl_141;
  wire and_dcpl_142;
  wire and_dcpl_143;
  wire and_dcpl_145;
  wire and_dcpl_146;
  wire and_dcpl_148;
  wire and_dcpl_150;
  wire and_dcpl_152;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire and_dcpl_159;
  wire and_dcpl_162;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_166;
  wire and_dcpl_167;
  wire and_dcpl_169;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire or_tmp;
  wire and_dcpl_172;
  wire or_tmp_12;
  wire mux_tmp_6;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_195;
  wire and_dcpl_213;
  wire or_dcpl_309;
  wire and_dcpl_215;
  wire and_dcpl_217;
  wire and_dcpl_249;
  wire and_dcpl_283;
  wire or_tmp_21;
  wire mux_tmp_7;
  wire and_dcpl_292;
  wire and_dcpl_293;
  wire and_dcpl_295;
  wire and_dcpl_296;
  wire and_dcpl_298;
  wire and_dcpl_300;
  wire and_dcpl_305;
  wire and_dcpl_317;
  wire and_dcpl_320;
  wire and_dcpl_342;
  wire and_dcpl_343;
  wire and_dcpl_346;
  wire and_dcpl_354;
  wire and_dcpl_360;
  wire and_dcpl_362;
  wire and_dcpl_365;
  wire and_dcpl_367;
  wire and_dcpl_369;
  wire and_dcpl_376;
  wire and_dcpl_377;
  wire and_dcpl_409;
  wire and_dcpl_418;
  wire and_dcpl_424;
  wire and_dcpl_427;
  wire and_dcpl_440;
  wire and_dcpl_443;
  wire and_dcpl_482;
  wire and_dcpl_492;
  wire and_dcpl_504;
  wire and_dcpl_509;
  wire and_dcpl_519;
  wire and_dcpl_541;
  wire and_dcpl_544;
  wire and_dcpl_554;
  wire and_dcpl_557;
  wire and_dcpl_564;
  wire and_dcpl_567;
  wire and_dcpl_581;
  wire or_tmp_35;
  wire or_tmp_40;
  wire mux_tmp_17;
  wire or_tmp_45;
  wire or_tmp_50;
  wire mux_tmp_20;
  wire or_tmp_56;
  wire or_tmp_57;
  wire or_tmp_60;
  wire mux_tmp_25;
  wire mux_tmp_26;
  wire or_tmp_85;
  wire or_tmp_87;
  wire or_dcpl_471;
  wire or_dcpl_475;
  wire or_dcpl_477;
  wire or_dcpl_480;
  wire or_dcpl_481;
  wire or_dcpl_483;
  wire or_dcpl_485;
  wire or_dcpl_489;
  wire or_dcpl_582;
  wire or_dcpl_587;
  wire or_dcpl_679;
  wire or_dcpl_684;
  wire and_dcpl_634;
  wire or_dcpl_694;
  wire or_tmp_89;
  wire or_tmp_90;
  wire or_tmp_91;
  wire or_tmp_92;
  wire or_tmp_95;
  wire or_tmp_96;
  wire mux_tmp_83;
  wire or_tmp_99;
  wire mux_tmp_85;
  wire mux_tmp_89;
  wire mux_tmp_99;
  wire nor_tmp_17;
  wire or_tmp_116;
  wire mux_tmp_139;
  wire mux_tmp_140;
  wire nor_tmp_19;
  wire mux_tmp_142;
  wire mux_tmp_143;
  wire or_tmp_129;
  wire mux_tmp_147;
  wire mux_tmp_150;
  wire mux_tmp_151;
  wire mux_tmp_152;
  wire mux_tmp_156;
  wire mux_tmp_161;
  wire not_tmp_277;
  wire or_tmp_147;
  wire nor_tmp_31;
  wire not_tmp_279;
  wire or_tmp_159;
  wire or_tmp_165;
  wire not_tmp_286;
  wire or_dcpl_700;
  wire or_dcpl_708;
  wire and_dcpl_750;
  wire or_dcpl_718;
  wire and_dcpl_832;
  wire and_dcpl_875;
  wire out_adp_set_value_ac_float_mux_95_tmp_3;
  wire out_adp_set_value_ac_float_mux_94_tmp_3;
  wire out_adp_set_value_ac_float_mux_93_tmp_3;
  wire out_adp_set_value_ac_float_mux_92_tmp_3;
  wire out_adp_set_value_ac_float_mux_91_tmp_3;
  wire out_adp_set_value_ac_float_mux_90_tmp_3;
  wire out_adp_set_value_ac_float_mux_89_tmp_3;
  wire out_adp_set_value_ac_float_mux_88_tmp_3;
  wire out_adp_set_value_ac_float_mux_87_tmp_3;
  wire out_adp_set_value_ac_float_mux_86_tmp_3;
  wire out_adp_set_value_ac_float_mux_85_tmp_3;
  wire out_adp_set_value_ac_float_mux_84_tmp_3;
  wire out_adp_set_value_ac_float_mux_83_tmp_3;
  wire out_adp_set_value_ac_float_mux_82_tmp_3;
  wire out_adp_set_value_ac_float_mux_81_tmp_3;
  wire out_adp_set_value_ac_float_mux_80_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_95_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_94_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_93_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_92_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_91_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_90_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_89_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_88_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_87_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_86_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_85_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_84_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_83_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_82_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_81_tmp_3;
  wire out_adp_set_value_ac_float_1_mux_80_tmp_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_1;
  reg NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2;
  wire NMP_UpdateFSM_case_11_time_end_lpi_1_dfm_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_1;
  reg NMP_UpdateFSM_switch_lp_equal_tmp_1;
  reg NMP_UpdateFSM_switch_lp_equal_tmp_1_1;
  reg NMP_UpdateFSM_switch_lp_equal_tmp_4_1;
  reg NMP_UpdateFSM_switch_lp_or_tmp_1;
  reg NMP_UpdateFSM_switch_lp_nor_tmp_1;
  reg NMP_UpdateFSM_switch_lp_equal_tmp_2_1;
  reg NMP_UpdateFSM_switch_lp_equal_tmp_3_1;
  reg NMP_UpdateFSM_switch_lp_equal_tmp_5_1;
  reg NMP_UpdateFSM_switch_lp_equal_tmp_6_1;
  reg next_state_3_lpi_1_dfm_3;
  reg nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1;
  reg ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_12;
  reg ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_12;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_16_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_15_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_14_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_14_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_13_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_13_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_12_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_11_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_10_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_9_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_9_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_8_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_7_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_7_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_6_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_5_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_4_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_4_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_3_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_3_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_2_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_2_itm_1;
  wire [3:0] out_adp_set_value_ac_float_exp_tmp_1_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_16_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_15_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_15_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_14_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_13_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_13_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_12_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_12_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_11_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_11_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_10_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_9_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_9_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_8_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_7_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_7_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_6_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_5_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_5_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_4_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_3_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_2_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1;
  wire [3:0] out_adp_set_value_ac_float_1_exp_tmp_1_lpi_1_dfm_4_1_mx0;
  reg in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_18;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_18;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_18;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_18;
  reg NMP_RunFSM_switch_lp_or_tmp_17;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_18;
  wire NMP_UpdateFSM_switch_lp_equal_tmp_7;
  wire NMP_UpdateFSM_switch_lp_equal_tmp_8;
  wire NMP_UpdateFSM_switch_lp_equal_tmp_10;
  wire NMP_UpdateFSM_switch_lp_equal_tmp_11;
  wire NMP_UpdateFSM_switch_lp_equal_tmp_9;
  wire NMP_UpdateFSM_switch_lp_equal_tmp_12;
  wire NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_6_cse_1;
  wire NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_7_cse_1;
  wire NMP_UpdateFSM_switch_lp_equal_tmp_13;
  wire NMP_RunFSM_switch_lp_equal_tmp_15;
  wire NMP_RunFSM_switch_lp_equal_tmp_14;
  wire NMP_RunFSM_switch_lp_equal_tmp_16;
  wire state_3_sva_mx1;
  wire state_1_sva_mx1;
  wire state_2_sva_mx1;
  wire state_0_sva_mx1;
  wire NMP_RunFSM_switch_lp_equal_tmp_22;
  wire NMP_RunFSM_switch_lp_equal_tmp_18_1;
  wire NMP_RunFSM_switch_lp_equal_tmp_20;
  wire NMP_RunFSM_switch_lp_equal_tmp_23;
  wire NMP_RunFSM_switch_lp_equal_tmp_17;
  wire NMP_RunFSM_switch_lp_equal_tmp_19;
  wire NMP_RunFSM_switch_lp_equal_tmp_21;
  wire NMP_RunFSM_switch_lp_equal_tmp_24;
  wire NMP_RunFSM_switch_lp_equal_tmp_25;
  wire NMP_RunFSM_switch_lp_or_tmp_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_1;
  wire NMP_ComputeSoftmaxMax_for_if_slc_NMP_ComputeSoftmaxMax_for_16_acc_1_27_svs_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_4;
  wire max_value_26_0_sva_dfm_14_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_14_25_0_mx0;
  reg max_value_26_0_sva_dfm_13_1_26;
  reg [25:0] max_value_26_0_sva_dfm_13_1_25_0;
  reg [26:0] NMP_ComputeSoftmaxMax_for_asn_13_itm_3;
  wire out_float_round_32_rnd_ovfl_sva_1;
  wire out_float_round_32_rnd_ovfl_15_sva_1;
  wire out_float_round_32_rnd_ovfl_14_sva_1;
  wire out_float_round_32_rnd_ovfl_13_sva_1;
  wire out_float_round_32_rnd_ovfl_12_sva_1;
  wire out_float_round_32_rnd_ovfl_11_sva_1;
  wire out_float_round_32_rnd_ovfl_10_sva_1;
  wire out_float_round_32_rnd_ovfl_9_sva_1;
  wire out_float_round_32_rnd_ovfl_8_sva_1;
  wire out_float_round_32_rnd_ovfl_7_sva_1;
  wire out_float_round_32_rnd_ovfl_6_sva_1;
  wire out_float_round_32_rnd_ovfl_5_sva_1;
  wire out_float_round_32_rnd_ovfl_4_sva_1;
  wire out_float_round_32_rnd_ovfl_3_sva_1;
  wire out_float_round_32_rnd_ovfl_2_sva_1;
  wire out_float_round_32_rnd_ovfl_1_sva_1;
  wire out_float_round_32_1_rnd_ovfl_sva_1;
  wire out_float_round_32_1_rnd_ovfl_15_sva_1;
  wire out_float_round_32_1_rnd_ovfl_14_sva_1;
  wire out_float_round_32_1_rnd_ovfl_13_sva_1;
  wire out_float_round_32_1_rnd_ovfl_12_sva_1;
  wire out_float_round_32_1_rnd_ovfl_11_sva_1;
  wire out_float_round_32_1_rnd_ovfl_10_sva_1;
  wire out_float_round_32_1_rnd_ovfl_9_sva_1;
  wire out_float_round_32_1_rnd_ovfl_8_sva_1;
  wire out_float_round_32_1_rnd_ovfl_7_sva_1;
  wire out_float_round_32_1_rnd_ovfl_6_sva_1;
  wire out_float_round_32_1_rnd_ovfl_5_sva_1;
  wire out_float_round_32_1_rnd_ovfl_4_sva_1;
  wire out_float_round_32_1_rnd_ovfl_3_sva_1;
  wire out_float_round_32_1_rnd_ovfl_2_sva_1;
  wire out_float_round_32_1_rnd_ovfl_1_sva_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_17_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_17;
  reg NMP_RunFSM_switch_lp_or_tmp_16;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17;
  wire max_value_26_0_sva_dfm_12_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_12_25_0_mx0;
  wire max_value_26_0_sva_dfm_11_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_11_25_0_mx0;
  wire max_value_26_0_sva_dfm_10_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_10_25_0_mx0;
  reg [33:0] NMP_ComputeSoftmaxSum_for_acc_7_itm_1;
  wire [35:0] nl_NMP_ComputeSoftmaxSum_for_acc_7_itm_1;
  reg [33:0] NMP_ComputeSoftmaxSum_for_acc_8_itm_1;
  wire [35:0] nl_NMP_ComputeSoftmaxSum_for_acc_8_itm_1;
  reg [33:0] NMP_ComputeSoftmaxSum_for_acc_9_itm_1;
  wire [35:0] nl_NMP_ComputeSoftmaxSum_for_acc_9_itm_1;
  reg [33:0] NMP_ComputeSoftmaxSum_for_acc_11_itm_1;
  wire [35:0] nl_NMP_ComputeSoftmaxSum_for_acc_11_itm_1;
  reg [32:0] NMP_ComputeSoftmaxSum_for_acc_12_itm_1;
  wire [33:0] nl_NMP_ComputeSoftmaxSum_for_acc_12_itm_1;
  reg [32:0] NMP_ComputeSoftmaxSum_for_acc_13_itm_1;
  wire [33:0] nl_NMP_ComputeSoftmaxSum_for_acc_13_itm_1;
  wire [2:0] nmp_config_mode_sva_mx1;
  wire max_value_26_0_sva_dfm_8_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_8_25_0_mx0;
  wire max_value_26_0_sva_dfm_7_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_7_25_0_mx0;
  reg max_value_26_0_sva_dfm_6_1_26;
  reg [25:0] max_value_26_0_sva_dfm_6_1_25_0;
  wire max_value_26_0_sva_dfm_5_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_5_25_0_mx0;
  reg [26:0] input_fixed_6_26_0_sva;
  wire max_value_26_0_sva_dfm_4_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_4_25_0_mx0;
  reg [26:0] input_fixed_5_26_0_sva;
  wire max_value_26_0_sva_dfm_3_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_3_25_0_mx0;
  reg [26:0] input_fixed_4_26_0_sva;
  wire [25:0] max_value_26_0_sva_dfm_1_25_0_mx0;
  reg [26:0] input_fixed_2_26_0_sva;
  wire NMP_ComputeSoftmaxMax_for_if_less_14_ssc_1;
  reg [26:0] input_fixed_0_26_0_sva;
  reg state_2_sva;
  reg state_1_sva;
  reg state_3_sva;
  reg state_0_sva;
  wire [35:0] sum_exp_39_4_sva_1;
  wire [38:0] nl_sum_exp_39_4_sva_1;
  wire NMP_RunFSM_switch_lp_equal_tmp_13;
  reg NMP_RunFSM_switch_lp_conc_itm_16_3;
  reg NMP_RunFSM_switch_lp_conc_itm_16_2;
  reg NMP_RunFSM_switch_lp_conc_itm_16_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_15;
  reg NMP_RunFSM_switch_lp_conc_itm_16_0;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_15;
  reg while_while_nor_itm_16;
  reg while_stage_0_18;
  reg NMP_RunFSM_switch_lp_conc_itm_15_3;
  reg NMP_RunFSM_switch_lp_conc_itm_15_1;
  reg NMP_RunFSM_switch_lp_conc_itm_15_2;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_15;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_14;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_13;
  reg NMP_RunFSM_switch_lp_conc_itm_12_0;
  reg NMP_RunFSM_switch_lp_conc_itm_12_3;
  reg NMP_RunFSM_switch_lp_conc_itm_12_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_12;
  reg ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_4;
  reg NMP_RunFSM_switch_lp_conc_itm_12_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_12;
  reg [35:0] sum_exp_39_4_sva_st_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_11;
  reg while_stage_0_14;
  reg NMP_RunFSM_switch_lp_conc_itm_11_0;
  reg NMP_RunFSM_switch_lp_conc_itm_11_3;
  reg NMP_RunFSM_switch_lp_conc_itm_11_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11;
  reg NMP_RunFSM_switch_lp_conc_itm_11_2;
  reg NMP_RunFSM_switch_lp_conc_itm_10_0;
  reg NMP_RunFSM_switch_lp_conc_itm_10_1;
  reg NMP_RunFSM_switch_lp_conc_itm_10_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10;
  reg NMP_RunFSM_switch_lp_conc_itm_10_2;
  reg NMP_RunFSM_switch_lp_conc_itm_9_0;
  reg NMP_RunFSM_switch_lp_conc_itm_9_1;
  reg NMP_RunFSM_switch_lp_conc_itm_9_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
  reg NMP_RunFSM_switch_lp_conc_itm_9_2;
  reg NMP_RunFSM_switch_lp_conc_itm_8_0;
  reg NMP_RunFSM_switch_lp_conc_itm_8_3;
  reg NMP_RunFSM_switch_lp_conc_itm_8_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  reg NMP_RunFSM_switch_lp_conc_itm_7_0;
  reg NMP_RunFSM_switch_lp_conc_itm_7_1;
  reg NMP_RunFSM_switch_lp_conc_itm_7_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  reg NMP_RunFSM_switch_lp_conc_itm_4_0;
  reg NMP_RunFSM_switch_lp_conc_itm_4_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  reg while_stage_0_3;
  reg state_1_sva_dfm_1;
  reg while_stage_0_17;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_14;
  reg NMP_RunFSM_switch_lp_conc_itm_7_2;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_3;
  reg ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_0_3_itm_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_3;
  reg NMP_RunFSM_switch_lp_conc_itm_4_1;
  reg NMP_RunFSM_switch_lp_conc_itm_4_2;
  reg NMP_RunFSM_switch_lp_conc_itm_3_0;
  reg NMP_RunFSM_switch_lp_conc_itm_3_3;
  reg while_while_nor_itm_15;
  reg NMP_RunFSM_switch_lp_conc_itm_8_2;
  reg NMP_RunFSM_switch_lp_conc_itm_6_3;
  reg NMP_RunFSM_switch_lp_conc_itm_6_0;
  reg NMP_RunFSM_switch_lp_conc_itm_6_2;
  reg NMP_RunFSM_switch_lp_conc_itm_6_1;
  reg NMP_RunFSM_switch_lp_conc_itm_15_0;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_10;
  reg ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_10;
  reg ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_2_1;
  reg [35:0] sum_exp_39_4_sva_st_2;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_2;
  reg ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_0_3_itm_2;
  reg NMP_RunFSM_switch_lp_conc_itm_3_2;
  reg while_while_nor_itm_14;
  reg while_stage_0_16;
  reg NMP_RunFSM_switch_lp_conc_itm_5_3;
  reg NMP_RunFSM_switch_lp_conc_itm_5_0;
  reg NMP_RunFSM_switch_lp_conc_itm_5_2;
  reg NMP_RunFSM_switch_lp_conc_itm_5_1;
  reg NMP_RunFSM_switch_lp_conc_itm_14_2;
  reg NMP_RunFSM_switch_lp_conc_itm_14_0;
  reg NMP_RunFSM_switch_lp_conc_itm_14_3;
  reg NMP_RunFSM_switch_lp_conc_itm_14_1;
  reg NMP_RunFSM_switch_lp_conc_itm_2_0;
  reg NMP_RunFSM_switch_lp_conc_itm_2_1;
  reg NMP_RunFSM_switch_lp_conc_itm_2_2;
  reg NMP_RunFSM_switch_lp_conc_itm_2_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_10;
  reg ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_9;
  reg while_stage_0_9;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1;
  wire [7:0] nl_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1;
  reg while_while_nor_itm_13;
  reg while_stage_0_15;
  reg NMP_RunFSM_switch_lp_conc_itm_13_2;
  reg NMP_RunFSM_switch_lp_conc_itm_13_0;
  reg NMP_RunFSM_switch_lp_conc_itm_13_3;
  reg NMP_RunFSM_switch_lp_conc_itm_13_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_8;
  reg NMP_RunFSM_switch_lp_conc_itm_3_1;
  reg while_while_nor_itm_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_2;
  reg while_stage_0_5;
  reg while_while_nor_itm_11;
  reg while_stage_0_13;
  reg while_while_nor_itm_10;
  reg while_stage_0_12;
  reg while_while_nor_itm_9;
  reg while_stage_0_11;
  reg while_while_nor_itm_8;
  reg while_stage_0_10;
  reg while_while_nor_itm_7;
  reg while_while_nor_itm_6;
  reg while_stage_0_8;
  reg while_while_nor_itm_5;
  reg while_stage_0_7;
  reg while_while_nor_itm_4;
  reg while_stage_0_6;
  reg while_while_nor_itm_3;
  reg while_while_nor_itm_2;
  reg while_stage_0_4;
  reg while_while_nor_itm_1;
  reg NMP_RunFSM_switch_lp_conc_itm_17_0;
  reg while_while_nor_itm_17;
  reg while_stage_0_19;
  reg while_while_and_itm_17;
  reg nmp_config_is_valid_sva;
  reg is_start_sva;
  reg NMP_RunFSM_switch_lp_conc_itm_17_2;
  reg NMP_RunFSM_switch_lp_conc_itm_17_1;
  reg NMP_RunFSM_switch_lp_conc_itm_17_3;
  reg while_stage_0_20;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_15;
  reg [39:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_3;
  reg [39:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_2;
  reg [35:0] sum_exp_39_4_sva_st_3;
  reg [39:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs;
  reg NMP_ComputeSoftmaxMax_for_if_less_5_itm_1;
  reg NMP_ComputeSoftmaxMax_for_if_less_12_itm_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_15_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_14_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_13_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_12_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_11_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_10_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_9_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_8_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_7_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_6_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_5_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_4_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_3_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_2_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_out_float_m_4_1_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_15_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_14_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_13_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_12_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_11_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_10_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_9_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_8_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_7_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_6_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_5_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_4_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_3_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_2_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_1_sva_1;
  wire max_value_26_0_sva_dfm_1_26_1;
  wire NMP_RunFSM_switch_lp_and_2_rgt;
  wire [39:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qelse_acc_sdt;
  wire [40:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qelse_acc_sdt;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_mx0_39;
  wire [38:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_mx0_38_0;
  wire xor_3_ssc;
  reg reg_NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo_ir_15_cse;
  reg reg_NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo_ir_15_cse;
  reg reg_NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo_ir_15_cse;
  reg reg_NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo_ir_15_cse;
  reg reg_done_Push_mioi_iswt0_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_large_rsp_PopNB_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_large_req_Push_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  reg [39:0] reg_NMP_ComputeRMSNormalize_for_1_mul_cmp_15_b_cse;
  reg [39:0] reg_NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_b_cse;
  wire large_req_reg_write_data_data_and_cse;
  wire write_data_data_and_16_cse;
  wire input_fixed_and_cse;
  wire state_and_cse;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_cse;
  wire nmp_config_num_vector_1_and_cse;
  wire operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
  wire operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_1_cse;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_2_cse;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_cse;
  wire or_503_cse;
  wire rva_out_reg_data_and_1_cse;
  wire [26:0] input_fixed_mux_7_cse;
  wire [26:0] input_fixed_mux_5_cse;
  wire [26:0] input_fixed_mux_3_cse;
  wire [26:0] input_fixed_mux_1_cse;
  wire [26:0] input_fixed_mux_25_cse;
  wire [26:0] input_fixed_mux_23_cse;
  wire [26:0] input_fixed_mux_21_cse;
  wire [26:0] input_fixed_mux_19_cse;
  wire [26:0] input_fixed_mux_17_cse;
  wire [26:0] input_fixed_mux_15_cse;
  wire [26:0] input_fixed_mux_13_cse;
  wire [26:0] input_fixed_mux_11_cse;
  wire [26:0] input_fixed_mux_9_cse;
  wire or_803_cse;
  wire nand_7_cse;
  wire and_899_cse;
  wire or_801_cse;
  wire NMP_RunFSM_switch_lp_and_8_cse_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_24_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_23_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_22_itm_1;
  wire mux_110_cse;
  wire while_and_142_rgt;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_cse;
  wire mux_105_cse_1;
  wire mux_107_cse;
  wire mux_131_cse;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_cse;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_1_cse;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_2_cse;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_3_cse;
  wire mux_49_cse;
  wire or_533_cse;
  wire [39:0] sum_exp_reciprocal_mux_rmff;
  wire [39:0] rms_reciprocal_mux_rmff;
  wire and_585_rmff;
  wire and_584_rmff;
  wire and_583_rmff;
  wire and_582_rmff;
  wire nor_206_rmff;
  wire and_591_rmff;
  wire and_590_rmff;
  wire and_588_rmff;
  wire and_587_rmff;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_17;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_17;
  reg large_req_reg_write_data_data_asn_itm_1;
  reg write_data_data_15_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_123_120_sva;
  wire [3:0] write_data_data_15_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_3_itm_1;
  reg write_data_data_14_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_115_112_sva;
  wire [3:0] write_data_data_14_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_6_itm_1;
  reg write_data_data_13_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_107_104_sva;
  wire [3:0] write_data_data_13_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_9_itm_1;
  reg write_data_data_12_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_99_96_sva;
  wire [3:0] write_data_data_12_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_12_itm_1;
  reg write_data_data_11_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_91_88_sva;
  wire [3:0] write_data_data_11_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_15_itm_1;
  reg write_data_data_10_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_83_80_sva;
  wire [3:0] write_data_data_10_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_18_itm_1;
  reg write_data_data_9_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_75_72_sva;
  wire [3:0] write_data_data_9_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_21_itm_1;
  reg write_data_data_8_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_67_64_sva;
  wire [3:0] write_data_data_8_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_24_itm_1;
  reg write_data_data_7_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_59_56_sva;
  wire [3:0] write_data_data_7_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_27_itm_1;
  reg write_data_data_6_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_51_48_sva;
  wire [3:0] write_data_data_6_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_30_itm_1;
  reg write_data_data_5_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_43_40_sva;
  wire [3:0] write_data_data_5_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_33_itm_1;
  reg write_data_data_4_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_35_32_sva;
  wire [3:0] write_data_data_4_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_36_itm_1;
  reg write_data_data_3_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_27_24_sva;
  wire [3:0] write_data_data_3_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_39_itm_1;
  reg write_data_data_2_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_19_16_sva;
  wire [3:0] write_data_data_2_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_42_itm_1;
  reg write_data_data_1_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_11_8_sva;
  wire [3:0] write_data_data_1_3_0_sva_dfm_1_mx1;
  reg large_req_reg_write_data_data_asn_45_itm_1;
  reg write_data_data_0_7_sva_dfm_1;
  reg [3:0] large_req_reg_write_data_data_3_0_sva;
  wire [3:0] write_data_data_0_3_0_sva_dfm_1_mx1;
  reg [1:0] large_req_reg_write_data_data_asn_1_itm_1_2_1;
  reg [1:0] write_data_data_15_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_1_itm_1_0;
  reg write_data_data_15_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_4_itm_1_2_1;
  reg [1:0] write_data_data_14_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_4_itm_1_0;
  reg write_data_data_14_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_7_itm_1_2_1;
  reg [1:0] write_data_data_13_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_7_itm_1_0;
  reg write_data_data_13_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_10_itm_1_2_1;
  reg [1:0] write_data_data_12_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_10_itm_1_0;
  reg write_data_data_12_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_13_itm_1_2_1;
  reg [1:0] write_data_data_11_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_13_itm_1_0;
  reg write_data_data_11_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_16_itm_1_2_1;
  reg [1:0] write_data_data_10_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_16_itm_1_0;
  reg write_data_data_10_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_19_itm_1_2_1;
  reg [1:0] write_data_data_9_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_19_itm_1_0;
  reg write_data_data_9_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_22_itm_1_2_1;
  reg [1:0] write_data_data_8_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_22_itm_1_0;
  reg write_data_data_8_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_25_itm_1_2_1;
  reg [1:0] write_data_data_7_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_25_itm_1_0;
  reg write_data_data_7_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_28_itm_1_2_1;
  reg [1:0] write_data_data_6_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_28_itm_1_0;
  reg write_data_data_6_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_31_itm_1_2_1;
  reg [1:0] write_data_data_5_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_31_itm_1_0;
  reg write_data_data_5_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_34_itm_1_2_1;
  reg [1:0] write_data_data_4_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_34_itm_1_0;
  reg write_data_data_4_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_37_itm_1_2_1;
  reg [1:0] write_data_data_3_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_37_itm_1_0;
  reg write_data_data_3_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_40_itm_1_2_1;
  reg [1:0] write_data_data_2_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_40_itm_1_0;
  reg write_data_data_2_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_43_itm_1_2_1;
  reg [1:0] write_data_data_1_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_43_itm_1_0;
  reg write_data_data_1_6_4_sva_dfm_1_0;
  reg [1:0] large_req_reg_write_data_data_asn_46_itm_1_2_1;
  reg [1:0] write_data_data_0_6_4_sva_dfm_1_2_1;
  reg large_req_reg_write_data_data_asn_46_itm_1_0;
  reg write_data_data_0_6_4_sva_dfm_1_0;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_45_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_43_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_41_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_39_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_37_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_35_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_33_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_31_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_29_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_27_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_25_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_23_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_21_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_19_itm_4;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_17_itm_4;
  reg [27:0] NMP_ComputeSoftmaxExp_for_1_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_1_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_16_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_16_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_15_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_15_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_14_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_14_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_13_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_13_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_12_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_12_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_11_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_11_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_10_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_10_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_9_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_9_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_8_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_8_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_7_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_7_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_6_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_6_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_5_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_5_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_4_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_4_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_3_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_3_acc_1_itm_1;
  reg [27:0] NMP_ComputeSoftmaxExp_for_2_acc_1_itm_1;
  wire [28:0] nl_NMP_ComputeSoftmaxExp_for_2_acc_1_itm_1;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_itm_11;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_60_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_58_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_56_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_54_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_52_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_50_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_48_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_46_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_44_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_42_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_40_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_38_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_36_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_34_itm_11;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_32_itm_11;
  reg [26:0] input_fixed_11_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_10_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_9_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_8_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_7_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_6_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_5_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_4_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_3_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_15_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_14_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_13_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_12_26_0_sva_dfm_2_1;
  reg [26:0] input_fixed_1_26_0_sva;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_17;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_17;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_17;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_17;
  reg rva_out_reg_data_0_sva_dfm_3_17;
  wire or_dcpl_742;
  reg NMP_RunFSM_switch_lp_equal_tmp_13_1;
  wire while_asn_736;
  reg NMP_RunFSM_switch_lp_equal_tmp_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_4;
  reg ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_4_39;
  reg [10:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_psp_sva;
  wire [11:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_psp_sva;
  wire [20:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_qif_ac_fixed_cctor_20_0_sva_1;
  wire [21:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_qif_ac_fixed_cctor_20_0_sva_1;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1_9_0;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_3;
  reg [10:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_itm;
  wire [11:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_itm;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TR000000;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_3;
  wire in_adp_is_zero_land_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_sva_1;
  wire in_adp_is_zero_land_15_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_15_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_15_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_15_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_15_sva_1;
  wire in_adp_is_zero_land_14_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_14_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_14_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_14_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_14_sva_1;
  wire in_adp_is_zero_land_13_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_13_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_13_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_13_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_13_sva_1;
  wire in_adp_is_zero_land_12_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_12_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_12_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_12_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_12_sva_1;
  wire in_adp_is_zero_land_11_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_11_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_11_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_11_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_11_sva_1;
  wire in_adp_is_zero_land_10_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_10_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_10_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_10_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_10_sva_1;
  wire in_adp_is_zero_land_9_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_9_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_9_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_9_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_9_sva_1;
  wire in_adp_is_zero_land_8_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_8_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_8_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_8_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_8_sva_1;
  wire in_adp_is_zero_land_7_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_7_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_7_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_7_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_7_sva_1;
  wire in_adp_is_zero_land_6_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_6_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_6_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_6_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_6_sva_1;
  wire in_adp_is_zero_land_5_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_5_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_5_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_5_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_5_sva_1;
  wire in_adp_is_zero_land_4_lpi_1_dfm_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_4_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_4_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_4_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_4_sva_1;
  reg [15:0] nmp_config_timestep_counter_sva;
  wire [39:0] operator_40_16_true_AC_TRN_AC_WRAP_rshift_itm;
  wire [39:0] operator_40_16_true_AC_TRN_AC_WRAP_1_rshift_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_itm;
  wire [26:0] NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_itm;
  wire [12:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_acc_itm;
  wire [13:0] nl_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_acc_itm;
  wire mux_216_itm;
  wire and_835_itm;
  wire [36:0] NMP_ComputeRMSSqrtRecip_variance_acc_itm;
  wire [37:0] nl_NMP_ComputeRMSSqrtRecip_variance_acc_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_16_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_15_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_14_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_13_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_12_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_11_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_10_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_9_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_8_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_7_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_6_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_5_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_4_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_3_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_2_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ComputeSoftmaxExp_for_1_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_16_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_15_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_14_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_13_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_12_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_11_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_10_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_9_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_8_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_7_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_6_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_5_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_4_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_3_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_2_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_for_1_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_16_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_15_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_14_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_13_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_12_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_11_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_10_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_9_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_8_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_7_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_6_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_5_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_4_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_3_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_2_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [31:0] NMP_ConvertOutputToAdpfloat_1_for_1_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [38:0] operator_40_0_false_AC_TRN_AC_WRAP_lshift_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_2_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_6_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_9_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_13_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_1_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_3_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_4_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_7_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_8_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_10_itm;
  wire NMP_ComputeSoftmaxMax_for_if_less_11_itm;
  wire and_dcpl_887;
  wire [7:0] z_out;
  wire [9:0] z_out_1;
  wire [38:0] z_out_2;
  wire and_dcpl_893;
  wire [5:0] rtn_out;
  reg [7:0] rva_out_reg_data_55_48_sva;
  reg [2:0] rva_out_reg_data_34_32_sva;
  reg [15:0] rva_out_reg_data_79_64_sva;
  reg [2:0] rva_out_reg_data_10_8_sva;
  reg rva_out_reg_data_0_sva;
  reg large_req_reg_write_data_data_63_sva;
  reg large_req_reg_write_data_data_71_sva;
  reg large_req_reg_write_data_data_55_sva;
  reg large_req_reg_write_data_data_79_sva;
  reg large_req_reg_write_data_data_47_sva;
  reg large_req_reg_write_data_data_87_sva;
  reg large_req_reg_write_data_data_39_sva;
  reg large_req_reg_write_data_data_95_sva;
  reg large_req_reg_write_data_data_31_sva;
  reg large_req_reg_write_data_data_103_sva;
  reg large_req_reg_write_data_data_23_sva;
  reg large_req_reg_write_data_data_111_sva;
  reg large_req_reg_write_data_data_15_sva;
  reg large_req_reg_write_data_data_119_sva;
  reg large_req_reg_write_data_data_7_sva;
  reg large_req_reg_write_data_data_127_sva;
  reg [2:0] nmp_config_mode_sva;
  reg [2:0] nmp_config_memory_index_1_sva;
  reg [7:0] nmp_config_num_vector_1_sva;
  reg [15:0] nmp_config_num_timestep_1_sva;
  reg [7:0] nmp_config_vector_counter_sva;
  reg [35:0] sum_sq_1_39_4_sva;
  reg [26:0] input_fixed_7_26_0_sva;
  reg [26:0] input_fixed_8_26_0_sva;
  reg [26:0] input_fixed_9_26_0_sva;
  reg [26:0] input_fixed_10_26_0_sva;
  reg [26:0] input_fixed_11_26_0_sva;
  reg [26:0] input_fixed_3_26_0_sva;
  reg [26:0] input_fixed_12_26_0_sva;
  reg [26:0] input_fixed_13_26_0_sva;
  reg [26:0] input_fixed_14_26_0_sva;
  reg [26:0] input_fixed_15_26_0_sva;
  reg [31:0] exp_values_7_sva;
  reg [31:0] exp_values_8_sva;
  reg [31:0] exp_values_6_sva;
  reg [31:0] exp_values_9_sva;
  reg [31:0] exp_values_5_sva;
  reg [31:0] exp_values_10_sva;
  reg [31:0] exp_values_4_sva;
  reg [31:0] exp_values_11_sva;
  reg [31:0] exp_values_3_sva;
  reg [31:0] exp_values_12_sva;
  reg [31:0] exp_values_2_sva;
  reg [31:0] exp_values_13_sva;
  reg [31:0] exp_values_1_sva;
  reg [31:0] exp_values_14_sva;
  reg [31:0] exp_values_0_sva;
  reg [31:0] exp_values_15_sva;
  reg NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs;
  reg next_state_1_lpi_1_dfm_3;
  reg [3:0] write_data_data_0_3_0_sva_dfm_1;
  reg [3:0] write_data_data_1_3_0_sva_dfm_1;
  reg [3:0] write_data_data_2_3_0_sva_dfm_1;
  reg [3:0] write_data_data_3_3_0_sva_dfm_1;
  reg [3:0] write_data_data_4_3_0_sva_dfm_1;
  reg [3:0] write_data_data_5_3_0_sva_dfm_1;
  reg [3:0] write_data_data_6_3_0_sva_dfm_1;
  reg [3:0] write_data_data_7_3_0_sva_dfm_1;
  reg [3:0] write_data_data_8_3_0_sva_dfm_1;
  reg [3:0] write_data_data_9_3_0_sva_dfm_1;
  reg [3:0] write_data_data_10_3_0_sva_dfm_1;
  reg [3:0] write_data_data_11_3_0_sva_dfm_1;
  reg [3:0] write_data_data_12_3_0_sva_dfm_1;
  reg [3:0] write_data_data_13_3_0_sva_dfm_1;
  reg [3:0] write_data_data_14_3_0_sva_dfm_1;
  reg [3:0] write_data_data_15_3_0_sva_dfm_1;
  reg [38:0] operator_40_0_false_AC_TRN_AC_WRAP_1_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_38_0_itm;
  reg [7:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_itm;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_itm;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_itm;
  reg ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_or_itm;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm;
  reg [7:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_itm;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_itm;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_itm;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm;
  reg [35:0] sum_exp_39_4_sva_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_14_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_15_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_16_1;
  reg NMP_RunFSM_switch_lp_or_tmp_1_1;
  reg NMP_RunFSM_switch_lp_or_tmp_2;
  reg NMP_RunFSM_switch_lp_or_tmp_3;
  reg NMP_RunFSM_switch_lp_or_tmp_4;
  reg NMP_RunFSM_switch_lp_or_tmp_5;
  reg NMP_RunFSM_switch_lp_or_tmp_6;
  reg NMP_RunFSM_switch_lp_or_tmp_7;
  reg NMP_RunFSM_switch_lp_or_tmp_8;
  reg NMP_RunFSM_switch_lp_or_tmp_9;
  reg NMP_RunFSM_switch_lp_or_tmp_10;
  reg NMP_RunFSM_switch_lp_or_tmp_11;
  reg NMP_RunFSM_switch_lp_or_tmp_12;
  reg NMP_RunFSM_switch_lp_or_tmp_13;
  reg NMP_RunFSM_switch_lp_or_tmp_14;
  reg NMP_RunFSM_switch_lp_or_tmp_15;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_15;
  reg NMP_RunFSM_switch_lp_equal_tmp_12_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_15;
  reg NMP_RunFSM_switch_lp_equal_tmp_11_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_15;
  reg NMP_RunFSM_switch_lp_equal_tmp_10_16;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_9_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_8_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_7_15;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_6_15;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_5_15;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_4_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_3_15;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_2_15;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_1;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_2;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_3;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_4;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_5;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_6;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_7;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_8;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_9;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_10;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_11;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_12;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_13;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_14;
  reg NMP_RunFSM_switch_lp_equal_tmp_1_15;
  reg [7:0] nmp_config_vector_counter_sva_3_1;
  wire [8:0] nl_nmp_config_vector_counter_sva_3_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_15_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_14_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_13_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_12_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_11_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_10_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_9_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_8_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_7_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_6_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_5_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_4_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_3_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_2_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_1_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_15_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_14_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_13_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_12_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_11_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_10_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_9_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_8_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_7_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_6_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_5_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_4_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_3_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_2_lpi_1_dfm_1_1;
  reg [3:0] NMP_ConvertOutputToAdpfloat_for_out_adp_man_1_lpi_1_dfm_1_1;
  reg [35:0] sum_sq_1_39_4_sva_2_1;
  reg [19:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_1_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_2_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_3_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_4_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_5_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_6_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_7_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_8_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_9_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_10_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_11_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_12_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_13_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_14_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_15_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeRMSNormalize_for_16_slc_55_24_ncse_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_1_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_2_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_3_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_4_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_5_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_6_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_7_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_8_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_9_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_10_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_11_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_12_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_13_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_14_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_15_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_1_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_2_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_3_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_4_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_5_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_6_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_7_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_8_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_9_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_10_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_11_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_12_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_13_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_14_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_15_slc_55_24_ncse_sva_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_16_slc_55_24_ncse_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_1_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_2_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_3_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_4_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_5_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_6_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_7_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_8_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_9_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_10_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_11_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_12_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_13_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_14_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_15_sva_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_sva_1;
  reg ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_1;
  reg ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_2;
  reg ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_3;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_2;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_3;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_4;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_5;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_6;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_7;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_8;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_9;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_10;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_11;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_12;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_13;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_14;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_15;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_3_16;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_2;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_3;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_4;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_5;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_6;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_7;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_8;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_9;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_10;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_11;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_12;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_13;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_14;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_15;
  reg [2:0] rva_out_reg_data_34_32_sva_dfm_3_16;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_2;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_3;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_4;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_5;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_6;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_7;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_8;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_9;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_10;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_11;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_12;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_13;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_14;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_15;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_3_16;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_2;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_3;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_4;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_5;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_6;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_7;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_8;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_9;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_10;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_11;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_12;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_13;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_14;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_15;
  reg [2:0] rva_out_reg_data_10_8_sva_dfm_3_16;
  reg rva_out_reg_data_0_sva_dfm_3_2;
  reg rva_out_reg_data_0_sva_dfm_3_3;
  reg rva_out_reg_data_0_sva_dfm_3_4;
  reg rva_out_reg_data_0_sva_dfm_3_5;
  reg rva_out_reg_data_0_sva_dfm_3_6;
  reg rva_out_reg_data_0_sva_dfm_3_7;
  reg rva_out_reg_data_0_sva_dfm_3_8;
  reg rva_out_reg_data_0_sva_dfm_3_9;
  reg rva_out_reg_data_0_sva_dfm_3_10;
  reg rva_out_reg_data_0_sva_dfm_3_11;
  reg rva_out_reg_data_0_sva_dfm_3_12;
  reg rva_out_reg_data_0_sva_dfm_3_13;
  reg rva_out_reg_data_0_sva_dfm_3_14;
  reg rva_out_reg_data_0_sva_dfm_3_15;
  reg rva_out_reg_data_0_sva_dfm_3_16;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_4;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_5;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_6;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_7;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_9;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_10;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_11;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_12;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_13;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_14;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_15;
  reg [1:0] NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_16;
  reg [7:0] NMP_PrepareReadReq_asn_1_itm_3;
  reg [15:0] NMP_PrepareReadReq_asn_2_itm_3;
  reg [15:0] NMP_PrepareReadReq_asn_2_itm_4;
  reg [9:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mux_1_itm_2;
  reg ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_itm_1;
  reg [5:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_6_1_itm_1;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_2;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_32_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_32_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_32_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_32_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_32_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_32_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_32_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_34_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_34_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_34_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_34_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_34_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_34_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_34_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_34_itm_10;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_36_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_36_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_36_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_36_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_36_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_36_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_36_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_38_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_38_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_38_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_38_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_38_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_38_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_38_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_40_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_40_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_40_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_40_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_40_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_40_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_40_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_42_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_42_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_42_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_42_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_42_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_42_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_42_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_44_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_44_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_44_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_44_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_44_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_44_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_44_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_46_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_46_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_46_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_46_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_46_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_46_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_46_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_48_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_48_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_48_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_48_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_48_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_48_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_48_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_50_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_50_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_50_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_50_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_50_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_50_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_50_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_52_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_52_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_52_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_52_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_52_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_52_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_52_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_54_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_54_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_54_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_54_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_54_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_54_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_54_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_56_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_56_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_56_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_56_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_56_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_56_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_56_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_58_itm_3;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_58_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_58_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_58_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_58_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_58_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_58_itm_9;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_60_itm_4;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_60_itm_5;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_60_itm_6;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_60_itm_7;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_60_itm_8;
  reg [26:0] NMP_ComputeRMSNormalize_for_asn_60_itm_9;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_1_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_2_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_3_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_4_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_5_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_6_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_7_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_8_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_9_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_10_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_11_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_12_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_13_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_14_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_15_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_itm_2;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_itm_3;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_2_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_16_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_16_itm_2;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_16_itm_3;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_6_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_7_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_17_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_17_itm_2;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_17_itm_3;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_18_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_18_itm_2;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_19_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_19_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_18_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_20_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_20_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_22_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_21_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_21_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_26_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_22_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_30_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_31_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_23_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_34_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_35_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_24_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_38_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_39_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_25_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_25_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_42_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_43_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_26_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_26_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_46_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_47_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_27_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_27_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_50_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_51_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_28_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_28_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_54_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_55_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_29_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_29_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_58_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_59_itm_1;
  reg [26:0] NMP_ComputeSoftmaxExp_for_asn_30_itm_2;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_62_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_63_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_8_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_9_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_7_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_6_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_11_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_5_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_12_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_4_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_13_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_3_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_14_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_2_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_15_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [8:0] NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000;
  reg [9:0] NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001;
  reg [8:0] NMP_ComputeSoftmaxExp_for_16_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1;
  reg [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_17_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_17_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_17_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_19_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_19_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_19_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_21_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_21_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_21_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_23_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_23_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_23_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_25_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_25_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_25_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_27_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_27_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_27_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_29_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_29_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_29_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_31_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_31_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_31_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_33_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_33_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_33_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_35_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_35_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_35_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_37_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_37_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_37_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_39_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_39_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_39_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_41_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_41_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_41_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_43_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_43_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_43_itm_3;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_45_itm_1;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_45_itm_2;
  reg [31:0] NMP_ComputeSoftmaxNormalize_for_asn_45_itm_3;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_1_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_2_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_3_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_4_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_5_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_6_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_7_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_8_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_9_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_10_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_11_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_12_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_13_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_14_itm_1;
  reg [4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_15_itm_1;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_2;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_3;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_4;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_5;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_6;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_7;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_9;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_10;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_11;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_12;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_13;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_14;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_15;
  reg [1:0] NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_16;
  reg [7:0] NMP_PrepareWriteReq_asn_1_itm_1;
  reg [7:0] NMP_PrepareWriteReq_asn_1_itm_2;
  reg [7:0] NMP_PrepareWriteReq_asn_1_itm_3;
  reg [7:0] NMP_PrepareWriteReq_asn_1_itm_4;
  reg [15:0] NMP_PrepareWriteReq_asn_2_itm_1;
  reg [15:0] NMP_PrepareWriteReq_asn_2_itm_2;
  reg [15:0] NMP_PrepareWriteReq_asn_2_itm_3;
  reg [15:0] NMP_PrepareWriteReq_asn_2_itm_4;
  reg [15:0] NMP_PrepareWriteReq_asn_2_itm_5;
  reg [15:0] NMP_PrepareWriteReq_asn_2_itm_6;
  reg [26:0] NMP_RunFSM_switch_lp_asn_104_itm_1;
  reg operator_3_false_operator_3_false_and_1_itm_1;
  reg operator_3_false_operator_3_false_and_1_itm_2;
  reg NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  reg [35:0] sum_exp_39_4_sva_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1;
  reg NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  reg while_while_and_itm_1;
  reg while_while_and_itm_2;
  reg while_while_and_itm_3;
  reg while_while_and_itm_4;
  reg while_while_and_itm_5;
  reg while_while_and_itm_6;
  reg while_while_and_itm_7;
  reg while_while_and_itm_8;
  reg while_while_and_itm_9;
  reg while_while_and_itm_10;
  reg while_while_and_itm_11;
  reg while_while_and_itm_12;
  reg while_while_and_itm_13;
  reg while_while_and_itm_14;
  reg while_while_and_itm_15;
  reg while_while_and_itm_16;
  reg [1:0] large_req_reg_write_data_data_62_60_sva_2_1;
  reg large_req_reg_write_data_data_62_60_sva_0;
  reg [1:0] large_req_reg_write_data_data_70_68_sva_2_1;
  reg large_req_reg_write_data_data_70_68_sva_0;
  reg [1:0] large_req_reg_write_data_data_54_52_sva_2_1;
  reg large_req_reg_write_data_data_54_52_sva_0;
  reg [1:0] large_req_reg_write_data_data_78_76_sva_2_1;
  reg large_req_reg_write_data_data_78_76_sva_0;
  reg [1:0] large_req_reg_write_data_data_46_44_sva_2_1;
  reg large_req_reg_write_data_data_46_44_sva_0;
  reg [1:0] large_req_reg_write_data_data_86_84_sva_2_1;
  reg large_req_reg_write_data_data_86_84_sva_0;
  reg [1:0] large_req_reg_write_data_data_38_36_sva_2_1;
  reg large_req_reg_write_data_data_38_36_sva_0;
  reg [1:0] large_req_reg_write_data_data_94_92_sva_2_1;
  reg large_req_reg_write_data_data_94_92_sva_0;
  reg [1:0] large_req_reg_write_data_data_30_28_sva_2_1;
  reg large_req_reg_write_data_data_30_28_sva_0;
  reg [1:0] large_req_reg_write_data_data_102_100_sva_2_1;
  reg large_req_reg_write_data_data_102_100_sva_0;
  reg [1:0] large_req_reg_write_data_data_22_20_sva_2_1;
  reg large_req_reg_write_data_data_22_20_sva_0;
  reg [1:0] large_req_reg_write_data_data_110_108_sva_2_1;
  reg large_req_reg_write_data_data_110_108_sva_0;
  reg [1:0] large_req_reg_write_data_data_14_12_sva_2_1;
  reg large_req_reg_write_data_data_14_12_sva_0;
  reg [1:0] large_req_reg_write_data_data_118_116_sva_2_1;
  reg large_req_reg_write_data_data_118_116_sva_0;
  reg [1:0] large_req_reg_write_data_data_6_4_sva_2_1;
  reg large_req_reg_write_data_data_6_4_sva_0;
  reg [1:0] large_req_reg_write_data_data_126_124_sva_2_1;
  reg large_req_reg_write_data_data_126_124_sva_0;
  reg out_float_round_32_1_if_m_1_1_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_1_sva_1_3_0;
  reg out_float_round_32_if_m_1_1_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_1_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_17_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_17_sva_1_3_0;
  reg out_float_round_32_if_m_1_17_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_17_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_16_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_16_sva_1_3_0;
  reg out_float_round_32_if_m_1_16_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_16_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_15_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_15_sva_1_3_0;
  reg out_float_round_32_if_m_1_15_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_15_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_14_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_14_sva_1_3_0;
  reg out_float_round_32_if_m_1_14_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_14_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_13_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_13_sva_1_3_0;
  reg out_float_round_32_if_m_1_13_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_13_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_12_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_12_sva_1_3_0;
  reg out_float_round_32_if_m_1_12_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_12_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_11_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_11_sva_1_3_0;
  reg out_float_round_32_if_m_1_11_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_11_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_10_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_10_sva_1_3_0;
  reg out_float_round_32_if_m_1_10_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_10_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_9_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_9_sva_1_3_0;
  reg out_float_round_32_if_m_1_9_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_9_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_8_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_8_sva_1_3_0;
  reg out_float_round_32_if_m_1_8_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_8_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_7_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_7_sva_1_3_0;
  reg out_float_round_32_if_m_1_7_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_7_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_6_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_6_sva_1_3_0;
  reg out_float_round_32_if_m_1_6_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_6_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_5_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_5_sva_1_3_0;
  reg out_float_round_32_if_m_1_5_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_5_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_4_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_4_sva_1_3_0;
  reg out_float_round_32_if_m_1_4_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_4_sva_1_3_0;
  reg out_float_round_32_1_if_m_1_3_sva_1_6;
  reg [3:0] out_float_round_32_1_if_m_1_3_sva_1_3_0;
  reg out_float_round_32_if_m_1_3_sva_1_6;
  reg [3:0] out_float_round_32_if_m_1_3_sva_1_3_0;
  reg ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_1_39;
  reg ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_2_39;
  reg ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_3_39;
  reg [34:0] sum_exp_39_4_sva_3_34_0;
  reg max_value_26_0_sva_dfm_2_1_26;
  reg [25:0] max_value_26_0_sva_dfm_2_1_25_0;
  reg max_value_26_0_sva_dfm_9_1_26;
  reg [25:0] max_value_26_0_sva_dfm_9_1_25_0;
  wire [3:0] write_data_data_15_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_14_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_13_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_12_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_11_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_10_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_9_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_8_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_7_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_6_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_5_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_4_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_3_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_2_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_1_3_0_sva_dfm_1_mx0w0;
  wire [3:0] write_data_data_0_3_0_sva_dfm_1_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_905_mx0w0;
  wire [1:0] write_data_data_15_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_15_6_4_sva_dfm_1_0_mx0w0;
  wire [1:0] write_data_data_0_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_0_6_4_sva_dfm_1_0_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_860_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_902_mx0w0;
  wire [1:0] write_data_data_14_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_14_6_4_sva_dfm_1_0_mx0w0;
  wire [1:0] write_data_data_1_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_1_6_4_sva_dfm_1_0_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_863_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_899_mx0w0;
  wire [1:0] write_data_data_13_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_13_6_4_sva_dfm_1_0_mx0w0;
  wire [1:0] write_data_data_2_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_2_6_4_sva_dfm_1_0_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_866_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_896_mx0w0;
  wire [1:0] write_data_data_12_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_12_6_4_sva_dfm_1_0_mx0w0;
  wire [1:0] write_data_data_3_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_3_6_4_sva_dfm_1_0_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_869_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_893_mx0w0;
  wire [1:0] write_data_data_11_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_11_6_4_sva_dfm_1_0_mx0w0;
  wire [1:0] write_data_data_4_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_4_6_4_sva_dfm_1_0_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_872_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_890_mx0w0;
  wire [1:0] write_data_data_10_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_10_6_4_sva_dfm_1_0_mx0w0;
  wire [1:0] write_data_data_5_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_5_6_4_sva_dfm_1_0_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_875_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_887_mx0w0;
  wire [1:0] write_data_data_9_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_9_6_4_sva_dfm_1_0_mx0w0;
  wire [1:0] write_data_data_6_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_6_6_4_sva_dfm_1_0_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_878_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_884_mx0w0;
  wire [1:0] write_data_data_8_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_8_6_4_sva_dfm_1_0_mx0w0;
  wire [1:0] write_data_data_7_6_4_sva_dfm_1_2_1_mx0w0;
  wire write_data_data_7_6_4_sva_dfm_1_0_mx0w0;
  wire NMP_RunFSM_switch_lp_mux1h_881_mx0w0;
  wire [7:0] nmp_config_vector_counter_sva_mx0w0;
  wire [7:0] nmp_config_vector_counter_sva_mx1;
  wire NMP_UpdateFSM_switch_lp_or_tmp_1_1;
  wire NMP_UpdateFSM_switch_lp_nor_tmp_1_1;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_1_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_1_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_2_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_2_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_3_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_3_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_4_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_4_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_5_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_5_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_6_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_6_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_7_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_7_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_8_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_8_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_9_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_9_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_10_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_10_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_11_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_11_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_12_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_12_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_13_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_13_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_14_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_14_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_15_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_15_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_acc_sdt_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_acc_sdt_sva_1;
  wire NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_1_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_1_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_2_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_2_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_3_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_3_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_4_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_4_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_5_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_5_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_6_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_6_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_7_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_7_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_8_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_8_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_9_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_9_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_10_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_10_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_11_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_11_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_12_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_12_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_13_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_13_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_14_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_14_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_15_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_15_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [4:0] out_adp_set_value_ac_float_1_acc_sdt_sva_1;
  wire [5:0] nl_out_adp_set_value_ac_float_1_acc_sdt_sva_1;
  wire NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  wire [18:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_mx0w0;
  wire signed [19:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_mx0w0;
  wire NMP_RunFSM_switch_lp_and_25_ssc_1;
  wire max_value_26_0_sva_dfm_9_1_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_9_1_25_0_mx0;
  wire nmp_config_adpbias_1_sva_dfm_3_1_mx0c0;
  wire nmp_config_adpbias_1_sva_dfm_3_1_mx0c1;
  wire nmp_config_adpbias_1_sva_dfm_3_1_mx0c2;
  wire [31:0] exp_values_15_sva_mx1;
  wire [31:0] exp_values_14_sva_mx1;
  wire [31:0] exp_values_13_sva_mx1;
  wire [31:0] exp_values_12_sva_mx1;
  wire [31:0] exp_values_11_sva_mx1;
  wire [31:0] exp_values_10_sva_mx1;
  wire [31:0] exp_values_9_sva_mx1;
  wire [31:0] exp_values_8_sva_mx1;
  wire [31:0] exp_values_7_sva_mx1;
  wire [31:0] exp_values_6_sva_mx1;
  wire [31:0] exp_values_5_sva_mx1;
  wire [31:0] exp_values_4_sva_mx1;
  wire [31:0] exp_values_3_sva_mx1;
  wire [31:0] exp_values_2_sva_mx1;
  wire [31:0] exp_values_1_sva_mx1;
  wire [31:0] exp_values_0_sva_mx1;
  wire max_value_26_0_sva_dfm_2_1_26_mx0;
  wire [25:0] max_value_26_0_sva_dfm_2_1_25_0_mx0;
  wire [35:0] sum_sq_1_39_4_sva_mx1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_1_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_1_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_1_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_1_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_2_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_2_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_2_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_2_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_3_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_3_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_3_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_3_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_4_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_4_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_4_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_4_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_5_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_5_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_5_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_5_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_6_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_6_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_6_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_6_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_7_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_7_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_7_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_7_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_8_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_8_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_8_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_8_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_9_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_9_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_9_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_9_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_10_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_10_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_10_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_10_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_11_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_11_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_11_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_11_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_12_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_12_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_12_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_12_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_13_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_13_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_13_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_13_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_14_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_14_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_14_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_14_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_15_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_15_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_15_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_15_sva_1;
  wire [4:0] out_adp_set_value_ac_float_exp_tmp_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_exp_tmp_sva_2;
  wire [3:0] out_adp_set_value_ac_float_ac_int_cctor_4_1_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_sva_1;
  wire out_adp_set_value_ac_float_lor_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_15_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_14_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_13_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_12_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_11_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_10_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_9_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_8_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_7_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_6_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_5_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_4_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_3_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_2_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_lor_1_lpi_1_dfm_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_1_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_1_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_1_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_1_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_2_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_2_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_2_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_2_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_3_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_3_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_3_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_3_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_4_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_4_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_4_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_4_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_5_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_5_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_5_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_5_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_6_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_6_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_6_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_6_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_7_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_7_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_7_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_7_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_8_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_8_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_8_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_8_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_9_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_9_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_9_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_9_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_10_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_10_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_10_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_10_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_11_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_11_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_11_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_11_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_12_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_12_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_12_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_12_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_13_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_13_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_13_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_13_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_14_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_14_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_14_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_14_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_15_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_15_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_15_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_15_sva_1;
  wire [4:0] out_adp_set_value_ac_float_1_exp_tmp_sva_2;
  wire [5:0] nl_out_adp_set_value_ac_float_1_exp_tmp_sva_2;
  wire [3:0] out_adp_set_value_ac_float_1_ac_int_cctor_4_1_sva_1;
  wire [4:0] nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_sva_1;
  wire out_adp_set_value_ac_float_1_lor_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_15_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_14_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_13_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_12_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_11_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_10_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_9_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_8_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_7_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_6_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_5_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_4_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_3_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_2_lpi_1_dfm_1;
  wire out_adp_set_value_ac_float_1_lor_1_lpi_1_dfm_1;
  wire next_state_0_lpi_1_dfm_4;
  wire next_state_2_lpi_1_dfm_4;
  wire next_state_3_lpi_1_dfm_4;
  wire in_adp_is_zero_land_3_lpi_1_dfm_1;
  wire in_adp_is_zero_land_2_lpi_1_dfm_1;
  wire in_adp_is_zero_land_1_lpi_1_dfm_1;
  wire NMP_RunFSM_switch_lp_or_861_cse_1;
  wire [18:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire signed [19:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire nmp_config_ConfigRead_unequal_tmp_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_1_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_1_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_1_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_1_sva_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_2_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_2_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_2_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_2_sva_1;
  wire [4:0] in_adp_to_ac_float_if_1_ac_int_cctor_4_0_3_sva_1;
  wire [5:0] nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_3_sva_1;
  wire [3:0] in_adp_to_ac_float_acc_sdt_3_sva_1;
  wire [4:0] nl_in_adp_to_ac_float_acc_sdt_3_sva_1;
  wire next_state_1_lpi_1_dfm_4;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_1_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_15_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_2_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_14_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_3_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_13_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_4_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_12_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_5_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_11_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_6_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_10_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_7_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_sva_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_8_sva_1;
  wire [25:0] NMP_ComputeSoftmaxMax_for_NMP_ComputeSoftmaxMax_for_and_psp_1;
  wire while_asn_728;
  wire while_asn_730;
  wire while_asn_732;
  wire while_asn_734;
  wire while_asn_738;
  wire while_asn_740;
  reg max_value_26_0_sva_26;
  reg [25:0] max_value_26_0_sva_25_0;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_9_0;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_10_5_0;
  wire NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_out_3;
  wire NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_out_2;
  wire [4:0] NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_out_3;
  wire [5:0] leading_sign_40_0_out_1;
  wire nmp_config_adpbias_1_and_ssc;
  reg reg_nmp_config_adpbias_1_ftd;
  reg [1:0] reg_nmp_config_adpbias_1_ftd_1;
  wire nmp_config_adpbias_1_sva_mx1_2;
  wire [1:0] nmp_config_adpbias_1_sva_mx1_1_0;
  wire nmp_config_adpbias_1_and_1_ssc;
  reg nmp_config_adpbias_1_sva_dfm_3_1_2;
  reg [1:0] nmp_config_adpbias_1_sva_dfm_3_1_1_0;
  wire [6:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_qif_acc_cse;
  wire [7:0] nl_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_qif_acc_cse;
  wire NMP_PrepareWriteReq_and_8_cse;
  wire NMP_PrepareWriteReq_and_9_cse;
  wire NMP_PrepareWriteReq_and_10_cse;
  wire NMP_PrepareWriteReq_and_11_cse;
  wire ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_7_cse;
  wire ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_5_cse;
  wire ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_6_cse;
  reg [26:0] reg_NMP_RunFSM_switch_lp_asn_104_itm_3_cse;
  wire NMP_ComputeRMSSqrtRecip_variance_and_1_ssc;
  reg [9:0] NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_36_27;
  reg [26:0] NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_26_0;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc;
  reg [3:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_12_9;
  reg [8:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_8_0;
  wire rva_out_reg_data_and_5_ssc;
  reg rva_out_reg_data_98_96_sva_dfm_3_1_2;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_1_1_0;
  wire NMP_PrepareReadReq_and_48_ssc;
  reg [1:0] NMP_PrepareReadReq_asn_1_itm_4_7_6;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_4_5_0;
  reg NMP_PrepareReadReq_asn_1_itm_7_7;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_11_5_0;
  reg [5:0] NMP_PrepareReadReq_asn_2_itm_5_15_10;
  reg [9:0] NMP_PrepareReadReq_asn_2_itm_5_9_0;
  wire NMP_PrepareReadReq_and_40_ssc;
  reg [6:0] NMP_PrepareReadReq_asn_2_itm_7_6_0;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc;
  reg [3:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_11_8;
  wire ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_29_ssc;
  reg ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_2;
  reg [1:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_1_0;
  wire ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_36_ssc;
  reg ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_14_itm_1_2;
  reg [1:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_14_itm_1_1_0;
  wire out_adp_set_value_ac_float_1_and_14_ssc;
  reg out_adp_set_value_ac_float_1_asn_15_itm_1_2;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_1_1_0;
  wire NMP_PrepareWriteReq_and_45_ssc;
  reg [1:0] NMP_PrepareWriteReq_asn_1_itm_5_7_6;
  reg [5:0] NMP_PrepareWriteReq_asn_1_itm_5_5_0;
  reg NMP_PrepareWriteReq_asn_1_itm_7_7;
  reg [8:0] NMP_PrepareWriteReq_asn_2_itm_7_15_7;
  reg [6:0] NMP_PrepareWriteReq_asn_2_itm_7_6_0;
  reg ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_39;
  reg [38:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_38_0;
  reg [3:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_7;
  reg [6:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_6_0;
  reg [9:0] NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_2_36_27;
  reg [26:0] NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_2_26_0;
  reg rva_out_reg_data_98_96_sva_dfm_3_2_2;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_2_1_0;
  reg NMP_PrepareReadReq_asn_1_itm_8_7;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_12_5_0;
  reg [5:0] NMP_PrepareReadReq_asn_2_itm_6_15_10;
  reg [9:0] NMP_PrepareReadReq_asn_2_itm_6_9_0;
  reg [6:0] NMP_PrepareReadReq_asn_2_itm_8_6_0;
  reg [3:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_1_itm_1_12_9;
  reg [8:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_1_itm_1_8_0;
  reg [3:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_2_itm_1_10_7;
  reg [6:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_2_itm_1_6_0;
  wire out_adp_set_value_ac_float_1_and_13_ssc;
  reg out_adp_set_value_ac_float_1_asn_15_itm_2_2;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_2_1_0;
  wire out_adp_set_value_ac_float_1_and_8_ssc;
  reg out_adp_set_value_ac_float_1_asn_15_itm_8_2;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_8_1_0;
  reg [1:0] NMP_PrepareWriteReq_asn_1_itm_6_7_6;
  reg [5:0] NMP_PrepareWriteReq_asn_1_itm_6_5_0;
  reg NMP_PrepareWriteReq_asn_1_itm_8_7;
  reg [8:0] NMP_PrepareWriteReq_asn_2_itm_8_15_7;
  reg [6:0] NMP_PrepareWriteReq_asn_2_itm_8_6_0;
  reg [1:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_7_6;
  reg [5:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_5_0;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_13_rsp_1;
  reg [8:0] NMP_PrepareWriteReq_asn_2_itm_9_rsp_0;
  reg [6:0] NMP_PrepareWriteReq_asn_2_itm_9_rsp_1;
  reg NMP_PrepareWriteReq_asn_1_itm_9_rsp_0;
  reg out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_0;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_1;
  wire out_adp_set_value_ac_float_1_and_7_ssc;
  reg [6:0] NMP_PrepareReadReq_asn_2_itm_9_rsp_1;
  reg NMP_PrepareReadReq_asn_1_itm_9_rsp_0;
  reg [1:0] NMP_PrepareReadReq_asn_1_itm_6_rsp_0;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_6_rsp_1;
  reg out_adp_set_value_ac_float_1_asn_15_itm_3_rsp_0;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_3_rsp_1;
  wire out_adp_set_value_ac_float_1_and_12_ssc;
  reg out_adp_set_value_ac_float_asn_15_itm_3_rsp_0;
  reg [1:0] out_adp_set_value_ac_float_asn_15_itm_3_rsp_1;
  reg rva_out_reg_data_98_96_sva_dfm_3_3_rsp_0;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_3_rsp_1;
  reg [5:0] reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_1;
  wire NMP_PrepareWriteReq_and_30_ssc;
  reg [8:0] reg_NMP_PrepareWriteReq_asn_2_itm_10_ftd;
  reg [6:0] reg_NMP_PrepareWriteReq_asn_2_itm_10_ftd_1;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_10_ftd;
  reg reg_out_adp_set_value_ac_float_1_asn_15_itm_10_ftd;
  reg [1:0] reg_out_adp_set_value_ac_float_1_asn_15_itm_10_ftd_1;
  reg reg_out_adp_set_value_ac_float_asn_15_itm_10_ftd;
  reg [1:0] reg_out_adp_set_value_ac_float_asn_15_itm_10_ftd_1;
  wire NMP_PrepareReadReq_and_32_ssc;
  reg [6:0] reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_1;
  reg reg_NMP_PrepareReadReq_asn_1_itm_10_ftd;
  reg reg_NMP_PrepareReadReq_asn_1_itm_10_ftd_1;
  wire out_adp_set_value_ac_float_1_and_11_ssc;
  reg reg_out_adp_set_value_ac_float_1_asn_15_itm_4_ftd;
  reg [1:0] reg_out_adp_set_value_ac_float_1_asn_15_itm_4_ftd_1;
  reg reg_out_adp_set_value_ac_float_asn_15_itm_4_ftd;
  reg [1:0] reg_out_adp_set_value_ac_float_asn_15_itm_4_ftd_1;
  reg reg_rva_out_reg_data_98_96_sva_dfm_3_4_ftd;
  reg [1:0] reg_rva_out_reg_data_98_96_sva_dfm_3_4_ftd_1;
  reg [5:0] reg_NMP_PrepareReadReq_asn_2_itm_7_ftd;
  reg [2:0] reg_NMP_PrepareReadReq_asn_2_itm_7_ftd_1;
  wire NMP_PrepareReadReq_and_7_ssc;
  reg NMP_PrepareReadReq_asn_1_itm_7_6;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_7_5_0;
  wire NMP_PrepareWriteReq_and_4_ssc;
  wire NMP_PrepareWriteReq_and_5_ssc;
  wire NMP_PrepareWriteReq_and_6_ssc;
  wire NMP_PrepareWriteReq_and_7_ssc;
  reg NMP_PrepareWriteReq_asn_1_itm_7_6;
  reg [5:0] NMP_PrepareWriteReq_asn_1_itm_7_5_0;
  reg rva_out_reg_data_98_96_sva_dfm_3_5_2;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_5_1_0;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_15_5_0;
  wire NMP_PrepareReadReq_and_29_ssc;
  reg [6:0] NMP_PrepareReadReq_asn_2_itm_11_6_0;
  reg out_adp_set_value_ac_float_asn_15_itm_5_2;
  reg [1:0] out_adp_set_value_ac_float_asn_15_itm_5_1_0;
  reg out_adp_set_value_ac_float_asn_15_itm_11_2;
  reg [1:0] out_adp_set_value_ac_float_asn_15_itm_11_1_0;
  wire out_adp_set_value_ac_float_1_and_10_ssc;
  reg out_adp_set_value_ac_float_1_asn_15_itm_5_2;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_5_1_0;
  reg out_adp_set_value_ac_float_1_asn_15_itm_11_2;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_11_1_0;
  reg NMP_PrepareWriteReq_asn_1_itm_11_7;
  wire NMP_PrepareWriteReq_and_27_ssc;
  reg [8:0] NMP_PrepareWriteReq_asn_2_itm_11_15_7;
  reg [6:0] NMP_PrepareWriteReq_asn_2_itm_11_6_0;
  reg NMP_PrepareReadReq_asn_1_itm_11_7;
  reg NMP_PrepareReadReq_asn_1_itm_11_6;
  reg NMP_PrepareReadReq_asn_1_itm_8_6;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_8_5_0;
  reg [5:0] NMP_PrepareReadReq_asn_2_itm_8_15_10;
  reg [2:0] NMP_PrepareReadReq_asn_2_itm_8_9_7;
  reg NMP_PrepareWriteReq_asn_1_itm_8_6;
  reg [5:0] NMP_PrepareWriteReq_asn_1_itm_8_5_0;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse;
  wire NMP_RunFSM_switch_lp_and_cse;
  wire large_req_reg_write_data_data_and_64_cse;
  wire in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
  wire in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
  wire NMP_PrepareWriteReq_and_12_cse;
  wire NMP_RunFSM_switch_lp_and_39_cse;
  wire rva_out_reg_data_and_6_cse;
  wire while_and_144_cse;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_cse;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_cse;
  wire NMP_RunFSM_switch_lp_and_43_cse;
  wire NMP_RunFSM_switch_lp_and_47_cse;
  wire NMP_RunFSM_switch_lp_and_51_cse;
  wire NMP_RunFSM_switch_lp_and_55_cse;
  wire NMP_RunFSM_switch_lp_and_56_cse;
  wire NMP_RunFSM_switch_lp_and_60_cse;
  wire NMP_ComputeRMSNormalize_for_and_cse;
  wire NMP_ComputeSoftmaxNormalize_for_and_cse;
  wire NMP_RunFSM_switch_lp_and_64_cse;
  wire NMP_RunFSM_switch_lp_and_68_cse;
  wire NMP_RunFSM_switch_lp_and_72_cse;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_2_cse;
  wire NMP_RunFSM_switch_lp_and_76_cse;
  wire NMP_RunFSM_switch_lp_and_80_cse;
  wire NMP_RunFSM_switch_lp_and_84_cse;
  wire NMP_RunFSM_switch_lp_and_88_cse;
  wire NMP_ComputeSoftmaxExp_for_and_cse;
  wire NMP_RunFSM_switch_lp_and_92_cse;
  wire NMP_RunFSM_switch_lp_and_96_cse;
  wire NMP_RunFSM_switch_lp_and_100_cse;
  wire NMP_RunFSM_switch_lp_and_104_cse;
  wire input_fixed_and_16_cse;
  wire while_if_and_17_cse;
  wire NMP_UpdateFSM_switch_lp_and_4_cse;
  wire large_req_reg_write_data_data_and_112_cse;
  wire large_req_reg_write_data_data_and_114_cse;
  wire while_if_and_12_cse;
  wire max_value_and_1_cse;
  wire while_if_and_13_cse;
  wire NMP_ComputeSoftmaxExp_for_and_17_cse;
  wire NMP_ComputeSoftmaxExp_for_and_22_cse;
  wire NMP_ComputeSoftmaxExp_for_and_29_cse;
  wire while_if_and_2_cse;
  wire NMP_PrepareWriteReq_and_15_cse;
  wire NMP_ComputeSoftmaxNormalize_for_and_32_cse;
  wire NMP_ComputeRMSNormalize_for_and_32_cse;
  wire NMP_PrepareReadReq_and_17_cse;
  wire rva_out_reg_data_and_12_cse;
  wire NMP_RunFSM_switch_lp_and_129_cse;
  wire while_if_and_6_cse;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_2_cse;
  wire NMP_ComputeSoftmaxSum_for_and_cse;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_6_cse;
  wire max_value_and_3_cse;
  wire while_if_and_3_cse;
  wire NMP_PrepareWriteReq_and_18_cse;
  wire NMP_ComputeSoftmaxNormalize_for_and_48_cse;
  wire NMP_ComputeSoftmaxExp_for_and_32_cse;
  wire NMP_ComputeSoftmaxExp_for_and_40_cse;
  wire NMP_ComputeSoftmaxExp_for_and_44_cse;
  wire NMP_ComputeRMSNormalize_for_and_48_cse;
  wire NMP_PrepareReadReq_and_20_cse;
  wire rva_out_reg_data_and_18_cse;
  wire NMP_RunFSM_switch_lp_and_135_cse;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_6_cse;
  wire while_if_and_7_cse;
  wire while_if_and_14_cse;
  wire ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_9_cse;
  wire while_if_and_10_cse;
  wire max_value_and_5_cse;
  wire while_if_and_4_cse;
  wire NMP_PrepareWriteReq_and_21_cse;
  wire NMP_ComputeSoftmaxNormalize_for_and_64_cse;
  wire NMP_ComputeSoftmaxExp_for_and_47_cse;
  wire NMP_ComputeRMSNormalize_for_and_64_cse;
  wire NMP_PrepareReadReq_and_23_cse;
  wire rva_out_reg_data_and_24_cse;
  wire NMP_RunFSM_switch_lp_and_158_cse;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_7_cse;
  wire while_if_and_8_cse;
  wire while_if_and_15_cse;
  wire max_value_and_7_cse;
  wire NMP_PrepareWriteReq_and_24_cse;
  wire NMP_ComputeRMSNormalize_for_and_80_cse;
  wire NMP_PrepareReadReq_and_26_cse;
  wire rva_out_reg_data_and_30_cse;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_9_cse;
  wire while_if_and_9_cse;
  wire while_if_and_11_cse;
  wire NMP_ComputeRMSNormalize_for_and_96_cse;
  wire rva_out_reg_data_and_36_cse;
  wire NMP_ComputeRMSNormalize_for_and_112_cse;
  wire rva_out_reg_data_and_42_cse;
  wire NMP_ComputeRMSNormalize_for_and_128_cse;
  wire rva_out_reg_data_and_48_cse;
  wire NMP_ComputeRMSNormalize_for_and_143_cse;
  wire rva_out_reg_data_and_54_cse;
  wire rva_out_reg_data_and_60_cse;
  wire NMP_PrepareWriteReq_and_41_cse;
  wire rva_out_reg_data_and_66_cse;
  wire NMP_PrepareWriteReq_and_44_cse;
  wire rva_out_reg_data_and_72_cse;
  wire NMP_PrepareWriteReq_and_47_cse;
  wire NMP_PrepareReadReq_and_47_cse;
  wire rva_out_reg_data_and_78_cse;
  wire NMP_PrepareWriteReq_and_50_cse;
  wire NMP_PrepareReadReq_and_50_cse;
  wire rva_out_reg_data_and_84_cse;
  wire NMP_PrepareWriteReq_and_53_cse;
  wire rva_out_reg_data_and_90_cse;
  wire NMP_PrepareWriteReq_and_56_cse;
  wire rva_out_reg_data_and_96_cse;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_2_cse;
  wire NMP_PrepareWriteReq_and_35_cse;
  wire NMP_PrepareReadReq_and_36_cse;
  wire NMP_PrepareWriteReq_and_38_cse;
  wire NMP_PrepareReadReq_and_39_cse;
  wire NMP_PrepareReadReq_and_44_cse;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_16_rsp_1;
  reg [8:0] NMP_PrepareWriteReq_asn_2_itm_12_rsp_0;
  reg [6:0] NMP_PrepareWriteReq_asn_2_itm_12_rsp_1;
  reg NMP_PrepareWriteReq_asn_1_itm_12_rsp_0;
  reg out_adp_set_value_ac_float_1_asn_15_itm_12_rsp_0;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_12_rsp_1;
  wire out_adp_set_value_ac_float_1_and_4_ssc;
  reg out_adp_set_value_ac_float_asn_15_itm_12_rsp_0;
  reg [1:0] out_adp_set_value_ac_float_asn_15_itm_12_rsp_1;
  wire out_adp_set_value_ac_float_and_4_ssc;
  reg [6:0] NMP_PrepareReadReq_asn_2_itm_12_rsp_1;
  reg out_adp_set_value_ac_float_1_asn_15_itm_6_rsp_0;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_6_rsp_1;
  wire out_adp_set_value_ac_float_1_and_9_ssc;
  reg out_adp_set_value_ac_float_asn_15_itm_6_rsp_0;
  reg [1:0] out_adp_set_value_ac_float_asn_15_itm_6_rsp_1;
  reg rva_out_reg_data_98_96_sva_dfm_3_6_rsp_0;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_6_rsp_1;
  reg NMP_PrepareReadReq_asn_1_itm_12_7_6_rsp_0;
  reg NMP_PrepareReadReq_asn_1_itm_12_7_6_rsp_1;
  reg NMP_PrepareWriteReq_asn_1_itm_9_rsp_1_rsp_0;
  reg [5:0] NMP_PrepareWriteReq_asn_1_itm_9_rsp_1_rsp_1;
  reg [5:0] NMP_PrepareReadReq_asn_2_itm_9_rsp_0_rsp_0;
  reg [2:0] NMP_PrepareReadReq_asn_2_itm_9_rsp_0_rsp_1;
  reg NMP_PrepareReadReq_asn_1_itm_9_rsp_1_rsp_0;
  reg [5:0] NMP_PrepareReadReq_asn_1_itm_9_rsp_1_rsp_1;
  reg [8:0] reg_NMP_PrepareWriteReq_asn_2_itm_13_ftd;
  reg [6:0] reg_NMP_PrepareWriteReq_asn_2_itm_13_ftd_1;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd;
  wire out_adp_set_value_ac_float_1_and_3_ssc;
  reg reg_out_adp_set_value_ac_float_1_asn_15_itm_13_ftd;
  reg [1:0] reg_out_adp_set_value_ac_float_1_asn_15_itm_13_ftd_1;
  wire out_adp_set_value_ac_float_and_3_ssc;
  reg reg_out_adp_set_value_ac_float_asn_15_itm_13_ftd;
  reg [1:0] reg_out_adp_set_value_ac_float_asn_15_itm_13_ftd_1;
  reg [6:0] reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_1;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_10_1_ftd;
  reg [5:0] reg_NMP_PrepareWriteReq_asn_1_itm_10_1_ftd_1;
  reg [5:0] reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_2;
  reg [2:0] reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_3;
  reg reg_rva_out_reg_data_98_96_sva_dfm_3_7_ftd;
  reg [1:0] reg_rva_out_reg_data_98_96_sva_dfm_3_7_ftd_1;
  reg reg_NMP_PrepareReadReq_asn_1_itm_13_ftd;
  reg reg_NMP_PrepareReadReq_asn_1_itm_13_ftd_1;
  reg rva_out_reg_data_98_96_sva_dfm_3_8_2;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_8_1_0;
  reg [6:0] NMP_PrepareReadReq_asn_2_itm_14_6_0;
  wire out_adp_set_value_ac_float_and_2_ssc;
  reg out_adp_set_value_ac_float_asn_15_itm_14_2;
  reg [1:0] out_adp_set_value_ac_float_asn_15_itm_14_1_0;
  wire out_adp_set_value_ac_float_1_and_2_ssc;
  reg out_adp_set_value_ac_float_1_asn_15_itm_14_2;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_14_1_0;
  reg NMP_PrepareWriteReq_asn_1_itm_14_7;
  reg [8:0] NMP_PrepareWriteReq_asn_2_itm_14_15_7;
  reg [6:0] NMP_PrepareWriteReq_asn_2_itm_14_6_0;
  reg reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_1_1;
  reg reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_0;
  wire input_fixed_and_37_cse;
  reg out_adp_set_value_ac_float_asn_15_itm_15_rsp_0;
  reg [1:0] out_adp_set_value_ac_float_asn_15_itm_15_rsp_1;
  reg out_adp_set_value_ac_float_1_asn_15_itm_15_rsp_0;
  reg [1:0] out_adp_set_value_ac_float_1_asn_15_itm_15_rsp_1;
  reg [8:0] NMP_PrepareWriteReq_asn_2_itm_15_rsp_0;
  reg [6:0] NMP_PrepareWriteReq_asn_2_itm_15_rsp_1;
  reg NMP_PrepareWriteReq_asn_1_itm_15_rsp_0;
  reg [6:0] NMP_PrepareReadReq_asn_2_itm_15_rsp_1;
  reg rva_out_reg_data_98_96_sva_dfm_3_9_rsp_0;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_9_rsp_1;
  reg NMP_PrepareReadReq_asn_1_itm_15_7_6_rsp_0;
  reg NMP_PrepareReadReq_asn_1_itm_15_7_6_rsp_1;
  reg NMP_PrepareWriteReq_asn_1_itm_11_6_0_rsp_0;
  reg [5:0] NMP_PrepareWriteReq_asn_1_itm_11_6_0_rsp_1;
  reg [5:0] NMP_PrepareReadReq_asn_2_itm_11_15_7_rsp_0;
  reg [2:0] NMP_PrepareReadReq_asn_2_itm_11_15_7_rsp_1;
  reg [6:0] reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_1;
  reg reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd;
  reg [1:0] reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1;
  reg reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd;
  reg [1:0] reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1;
  reg [8:0] reg_NMP_PrepareWriteReq_asn_2_itm_16_ftd;
  reg [6:0] reg_NMP_PrepareWriteReq_asn_2_itm_16_ftd_1;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd;
  reg reg_rva_out_reg_data_98_96_sva_dfm_3_10_ftd;
  reg [1:0] reg_rva_out_reg_data_98_96_sva_dfm_3_10_ftd_1;
  reg reg_NMP_PrepareReadReq_asn_1_itm_16_ftd;
  reg reg_NMP_PrepareReadReq_asn_1_itm_16_ftd_1;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_12_1_ftd;
  reg [5:0] reg_NMP_PrepareWriteReq_asn_1_itm_12_1_ftd_1;
  reg [5:0] reg_NMP_PrepareReadReq_asn_2_itm_12_ftd;
  reg [2:0] reg_NMP_PrepareReadReq_asn_2_itm_12_ftd_1;
  reg rva_out_reg_data_98_96_sva_dfm_3_11_2;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_11_1_0;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd_1_6;
  reg [5:0] reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd_1_5_0;
  reg [5:0] reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_8_3;
  reg [2:0] reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_2_0;
  reg rva_out_reg_data_98_96_sva_dfm_3_12_rsp_0;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_12_rsp_1;
  reg NMP_PrepareWriteReq_asn_1_itm_14_6_0_rsp_0;
  reg [5:0] NMP_PrepareWriteReq_asn_1_itm_14_6_0_rsp_1;
  reg [5:0] NMP_PrepareReadReq_asn_2_itm_14_15_7_rsp_0;
  reg [2:0] NMP_PrepareReadReq_asn_2_itm_14_15_7_rsp_1;
  reg reg_rva_out_reg_data_98_96_sva_dfm_3_13_ftd;
  reg [1:0] reg_rva_out_reg_data_98_96_sva_dfm_3_13_ftd_1;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_15_1_ftd;
  reg [5:0] reg_NMP_PrepareWriteReq_asn_1_itm_15_1_ftd_1;
  reg [5:0] reg_NMP_PrepareReadReq_asn_2_itm_15_ftd;
  reg [2:0] reg_NMP_PrepareReadReq_asn_2_itm_15_ftd_1;
  reg rva_out_reg_data_98_96_sva_dfm_3_14_2;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_14_1_0;
  reg [5:0] reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_8_3;
  reg [2:0] reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_2_0;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd_1_6;
  reg [5:0] reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd_1_5_0;
  reg rva_out_reg_data_98_96_sva_dfm_3_15_rsp_0;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_15_rsp_1;
  reg reg_rva_out_reg_data_98_96_sva_dfm_3_16_ftd;
  reg [1:0] reg_rva_out_reg_data_98_96_sva_dfm_3_16_ftd_1;
  reg rva_out_reg_data_98_96_sva_dfm_3_17_2;
  reg [1:0] rva_out_reg_data_98_96_sva_dfm_3_17_1_0;
  wire or_928_cse;
  wire or_929_cse;
  wire or_534_cse;
  wire and_936_cse;
  wire and_983_cse;
  wire and_1011_cse;
  wire mux_cse;
  wire and_1067_cse;
  wire and_1094_cse;
  wire or_1057_cse;
  wire nor_58_cse;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_15_itm_1_enexo;
  reg reg_out_float_round_32_if_m_1_1_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_out_float_round_32_if_m_1_1_sva_1_3_0_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_15_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_1_sva_1_3_0_enexo;
  reg reg_out_float_round_32_1_if_m_1_1_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_if_m_1_17_sva_1_6_enexo;
  reg reg_out_float_round_32_if_m_1_17_sva_1_3_0_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_17_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_14_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_17_sva_1_3_0_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_13_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_out_float_round_32_if_m_1_16_sva_1_3_0_enexo;
  reg reg_out_float_round_32_if_m_1_16_sva_1_6_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_16_sva_1_3_0_enexo;
  reg reg_out_float_round_32_1_if_m_1_16_sva_1_6_enexo;
  reg reg_out_float_round_32_if_m_1_15_sva_1_6_enexo;
  reg reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_3;
  reg reg_out_float_round_32_if_m_1_15_sva_1_3_0_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_12_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_15_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_15_sva_1_3_0_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_out_float_round_32_if_m_1_14_sva_1_3_0_enexo;
  reg reg_out_float_round_32_if_m_1_14_sva_1_6_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_14_sva_1_3_0_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_11_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_14_sva_1_6_enexo;
  reg reg_out_float_round_32_if_m_1_13_sva_1_3_0_enexo;
  reg reg_out_float_round_32_if_m_1_13_sva_1_6_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_10_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_13_sva_1_6_enexo;
  reg reg_out_float_round_32_1_if_m_1_13_sva_1_3_0_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_out_float_round_32_if_m_1_12_sva_1_3_0_enexo;
  reg reg_out_float_round_32_if_m_1_12_sva_1_6_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_12_sva_1_3_0_enexo;
  reg reg_out_float_round_32_1_if_m_1_12_sva_1_6_enexo;
  reg reg_out_float_round_32_if_m_1_11_sva_1_3_0_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_7;
  reg reg_out_float_round_32_if_m_1_11_sva_1_6_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_8_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_11_sva_1_6_enexo;
  reg reg_out_float_round_32_1_if_m_1_11_sva_1_3_0_enexo;
  reg reg_out_float_round_32_if_m_1_10_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1_enexo;
  reg reg_out_float_round_32_if_m_1_10_sva_1_3_0_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_10_sva_1_3_0_enexo;
  reg reg_out_float_round_32_1_if_m_1_10_sva_1_6_enexo;
  reg reg_out_float_round_32_if_m_1_9_sva_1_3_0_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_6_itm_1_enexo;
  reg reg_out_float_round_32_if_m_1_9_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_6_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_9_sva_1_3_0_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_9_sva_1_6_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1_enexo;
  reg reg_out_float_round_32_if_m_1_8_sva_1_3_0_enexo;
  reg reg_out_float_round_32_if_m_1_8_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_8_sva_1_3_0_enexo;
  reg reg_out_float_round_32_1_if_m_1_8_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1_enexo;
  reg reg_out_float_round_32_if_m_1_7_sva_1_3_0_enexo;
  reg reg_out_float_round_32_if_m_1_7_sva_1_6_enexo;
  reg reg_out_float_round_32_1_if_m_1_7_sva_1_6_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_4_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_7_sva_1_3_0_enexo;
  reg reg_out_float_round_32_if_m_1_6_sva_1_3_0_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_3_itm_1_enexo;
  reg reg_out_float_round_32_if_m_1_6_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_6_sva_1_3_0_enexo;
  reg reg_out_float_round_32_1_if_m_1_6_sva_1_6_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_if_m_1_5_sva_1_6_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_2_itm_1_enexo;
  reg reg_out_float_round_32_if_m_1_5_sva_1_3_0_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_5_sva_1_3_0_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_5_sva_1_6_enexo;
  reg reg_out_float_round_32_if_m_1_4_sva_1_6_enexo;
  reg reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_14;
  reg reg_out_float_round_32_if_m_1_4_sva_1_3_0_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_4_sva_1_6_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_4_sva_1_3_0_enexo;
  reg reg_out_float_round_32_if_m_1_3_sva_1_6_enexo;
  reg reg_out_float_round_32_if_m_1_3_sva_1_3_0_enexo;
  reg reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_itm_1_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo;
  reg reg_NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo;
  reg reg_out_float_round_32_1_if_m_1_3_sva_1_3_0_enexo;
  reg reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1_enexo;
  reg reg_out_float_round_32_1_if_m_1_3_sva_1_6_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_15_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_15_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_15_1_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_16_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_16_enexo;
  reg reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_enexo;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_3_enexo;
  reg reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_2_enexo;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_2_enexo;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_2_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_60_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_58_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_56_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_54_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_52_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_50_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_48_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_46_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_44_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_42_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_40_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_38_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_36_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_34_itm_10_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_32_itm_10_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_itm_10_enexo;
  reg reg_sum_exp_39_4_sva_st_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_3_enexo;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_1_enexo;
  reg reg_sum_exp_39_4_sva_st_2_enexo;
  reg reg_sum_exp_39_4_sva_st_1_enexo;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo;
  reg reg_max_value_26_0_1_enexo;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_30_itm_2_enexo;
  reg reg_while_stage_0_7_enexo;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo;
  reg reg_max_value_26_0_enexo;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_1;
  reg reg_max_value_26_0_1_enexo_1;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_1;
  reg reg_while_stage_0_7_enexo_1;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_1;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_1;
  reg reg_max_value_26_0_enexo_1;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_2;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_2;
  reg reg_max_value_26_0_1_enexo_2;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_2;
  reg reg_while_stage_0_7_enexo_2;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_2;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_2;
  reg reg_max_value_26_0_enexo_2;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_3;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_3;
  reg reg_max_value_26_0_1_enexo_3;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_3;
  reg reg_while_stage_0_7_enexo_3;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_3;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_3;
  reg reg_max_value_26_0_enexo_3;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_4;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_4;
  reg reg_max_value_26_0_1_enexo_4;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_4;
  reg reg_while_stage_0_7_enexo_4;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_4;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_4;
  reg reg_max_value_26_0_enexo_4;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_5;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_5;
  reg reg_max_value_26_0_1_enexo_5;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_5;
  reg reg_while_stage_0_7_enexo_5;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_5;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_5;
  reg reg_max_value_26_0_enexo_5;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_6;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_2_enexo;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_6;
  reg reg_max_value_26_0_1_enexo_6;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_6;
  reg reg_while_stage_0_7_enexo_6;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_6;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_6;
  reg reg_max_value_26_0_enexo_6;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_7;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_7;
  reg reg_max_value_26_0_1_enexo_7;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_2_enexo;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_7;
  reg reg_while_stage_0_7_enexo_7;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_7;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_7;
  reg reg_max_value_26_0_enexo_7;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_8;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_2_enexo;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_8;
  reg reg_max_value_26_0_1_enexo_8;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_8;
  reg reg_while_stage_0_7_enexo_8;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_8;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_8;
  reg reg_max_value_26_0_enexo_8;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_9;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_9;
  reg reg_max_value_26_0_1_enexo_9;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_9;
  reg reg_while_stage_0_7_enexo_9;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_9;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_9;
  reg reg_max_value_26_0_enexo_9;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_2_enexo;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_10;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_10;
  reg reg_max_value_26_0_1_enexo_10;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_10;
  reg reg_while_stage_0_7_enexo_10;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_10;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_10;
  reg reg_max_value_26_0_enexo_10;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_11;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_2_enexo;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_11;
  reg reg_max_value_26_0_1_enexo_11;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_11;
  reg reg_while_stage_0_7_enexo_11;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_11;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_11;
  reg reg_max_value_26_0_enexo_11;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_12;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_12;
  reg reg_max_value_26_0_1_enexo_12;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_12;
  reg reg_while_stage_0_7_enexo_12;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_12;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_12;
  reg reg_max_value_26_0_enexo_12;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_3_enexo;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_13;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_13;
  reg reg_max_value_26_0_1_enexo_13;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_13;
  reg reg_while_stage_0_7_enexo_13;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_13;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_13;
  reg reg_max_value_26_0_enexo_13;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_14;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_14;
  reg reg_max_value_26_0_1_enexo_14;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_14;
  reg reg_while_stage_0_7_enexo_14;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_3_enexo;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_14;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_14;
  reg reg_max_value_26_0_enexo_14;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_15;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_15;
  reg reg_max_value_26_0_1_enexo_15;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_15;
  reg reg_while_stage_0_7_enexo_15;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_15;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_15;
  reg reg_max_value_26_0_enexo_15;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_itm_3_enexo;
  reg reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_enexo;
  reg reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo_2;
  reg reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo;
  reg reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_enexo;
  reg reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_16;
  reg reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_16;
  reg reg_max_value_26_0_1_enexo_16;
  reg reg_max_value_26_0_sva_dfm_13_1_26_enexo_16;
  reg reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_16;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_16;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_30_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo_1;
  reg reg_max_value_26_0_sva_dfm_9_1_25_0_enexo;
  reg reg_NMP_ComputeSoftmaxMax_for_if_less_5_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo_1;
  reg reg_max_value_26_0_sva_dfm_9_1_26_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo_1;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxSum_for_acc_7_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_2_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_2_enexo;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_60_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_58_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_56_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_54_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_52_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_50_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_48_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_46_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_44_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_42_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_40_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_38_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_36_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_34_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_32_itm_9_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_itm_9_enexo;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_15_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_15_enexo;
  reg reg_sum_exp_39_4_sva_2_enexo;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_5_1_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_5_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_1_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_1_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_1_enexo_1;
  reg reg_max_value_26_0_sva_dfm_6_1_25_0_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_1_enexo;
  reg reg_input_fixed_14_26_0_enexo;
  reg reg_input_fixed_13_26_0_enexo;
  reg reg_input_fixed_12_26_0_enexo;
  reg reg_input_fixed_11_26_0_enexo;
  reg reg_input_fixed_10_26_0_enexo;
  reg reg_input_fixed_9_26_0_enexo;
  reg reg_input_fixed_8_26_0_enexo;
  reg reg_input_fixed_7_26_0_enexo;
  reg reg_input_fixed_6_26_0_enexo;
  reg reg_input_fixed_5_26_0_enexo;
  reg reg_input_fixed_4_26_0_enexo;
  reg reg_input_fixed_3_26_0_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_1_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_itm_1_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_60_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_58_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_56_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_54_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_52_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_50_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_48_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_46_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_44_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_42_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_40_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_38_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_36_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_34_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_32_itm_8_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_itm_8_enexo;
  reg reg_NMP_PrepareReadReq_asn_1_itm_13_1_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_14_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_14_enexo;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_2_enexo;
  reg reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_1_enexo;
  reg reg_sum_exp_39_4_sva_st_1_enexo_1;
  reg reg_input_fixed_15_26_0_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_12_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_12_1_enexo;
  reg reg_exp_values_15_enexo;
  reg reg_exp_values_14_enexo;
  reg reg_exp_values_13_enexo;
  reg reg_exp_values_12_enexo;
  reg reg_exp_values_11_enexo;
  reg reg_exp_values_10_enexo;
  reg reg_exp_values_9_enexo;
  reg reg_exp_values_8_enexo;
  reg reg_exp_values_7_enexo;
  reg reg_exp_values_6_enexo;
  reg reg_exp_values_5_enexo;
  reg reg_exp_values_4_enexo;
  reg reg_exp_values_3_enexo;
  reg reg_exp_values_2_enexo;
  reg reg_exp_values_1_enexo;
  reg reg_exp_values_0_enexo;
  reg reg_input_fixed_2_26_0_enexo;
  reg reg_input_fixed_1_26_0_enexo;
  reg reg_input_fixed_0_26_0_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_60_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_58_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_56_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_54_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_52_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_50_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_48_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_46_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_44_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_42_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_40_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_38_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_36_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_34_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_32_itm_7_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_itm_7_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_12_1_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_13_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_13_enexo;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1_enexo;
  reg reg_input_fixed_1_26_0_enexo_1;
  reg reg_NMP_ComputeRMSNormalize_for_asn_60_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_58_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_56_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_54_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_52_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_50_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_48_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_46_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_44_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_42_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_40_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_38_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_36_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_34_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_32_itm_6_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_itm_6_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_12_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_12_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_60_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_58_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_56_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_54_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_52_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_50_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_48_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_46_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_44_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_42_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_40_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_38_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_36_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_34_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_32_itm_5_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_itm_5_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_11_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_11_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_9_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_9_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_9_2_enexo;
  reg reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_17;
  reg reg_NMP_ComputeRMSNormalize_for_asn_58_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_56_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_54_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_52_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_50_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_48_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_46_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_44_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_42_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_40_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_38_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_36_itm_3_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_34_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_32_itm_4_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_itm_4_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_9_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_9_1_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_10_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_10_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo_2;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo_2;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo_2;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo_2;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo_2;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_2_enexo_1;
  reg reg_NMP_ComputeRMSNormalize_for_asn_34_itm_3_enexo;
  reg reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_1_enexo;
  reg reg_NMP_ComputeRMSNormalize_for_asn_itm_3_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_9_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_9_enexo;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_2_enexo_1;
  reg reg_NMP_ComputeSoftmaxExp_for_asn_itm_2_enexo_1;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_8_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_8_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_7_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_7_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_5_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_6_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_6_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_4_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_5_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_5_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_3_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_3_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_3_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_4_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_4_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_2_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_2_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_2_enexo_1;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_2_enexo_1;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_3_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_1_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_3_2_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_3_2_enexo;
  reg reg_nmp_config_timestep_counter_enexo;
  reg reg_nmp_config_vector_counter_enexo;
  reg reg_rva_out_reg_data_79_64_enexo;
  reg reg_rva_out_reg_data_55_48_enexo;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_1;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_1;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_1;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_1;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_2;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_2;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_2;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_2;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_3;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_3;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_3;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_3;
  reg reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_4;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mux_1_itm_2_enexo;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1_enexo;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1_enexo_1;
  reg reg_NMP_PrepareReadReq_asn_1_itm_12_1_enexo;
  reg reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_enexo;
  reg reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_1_enexo_1;
  reg reg_NMP_PrepareReadReq_asn_1_itm_11_1_enexo;
  reg reg_NMP_PrepareReadReq_asn_1_itm_10_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_8_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_8_1_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_8_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_7_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_7_1_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_7_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_6_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_6_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_5_1_enexo_1;
  reg reg_NMP_PrepareReadReq_asn_2_itm_5_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_5_1_enexo_1;
  reg reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_2_enexo_1;
  reg reg_NMP_PrepareReadReq_asn_2_itm_4_enexo;
  reg reg_NMP_PrepareReadReq_asn_1_itm_15_1_enexo;
  reg reg_NMP_PrepareReadReq_asn_1_itm_14_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_11_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_11_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_11_2_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_11_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_11_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_10_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_10_1_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_10_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_8_2_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_8_enexo;
  reg reg_NMP_PrepareReadReq_asn_1_itm_8_2_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_7_2_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_7_enexo;
  reg reg_NMP_PrepareReadReq_asn_1_itm_7_2_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_14_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_14_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_14_2_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_14_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_14_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_13_enexo;
  reg reg_NMP_PrepareWriteReq_asn_2_itm_13_1_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_13_1_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_10_2_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_10_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_12_2_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_12_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_13_2_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_13_enexo;
  reg reg_NMP_PrepareReadReq_asn_2_itm_15_enexo;
  reg reg_NMP_PrepareWriteReq_asn_1_itm_15_2_enexo;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_16_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_16_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_17_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_17_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_18_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_18_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_19_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_19_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_20_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_20_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_21_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_21_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_22_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_22_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_23_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_23_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_24_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_24_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_25_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_25_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_26_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_26_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_27_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_27_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_28_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_28_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_29_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_29_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_30_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_30_enex5;
  wire NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_31_enex5;
  wire NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_31_enex5;
  wire NMP_PrepareReadReq_and_55_enex5;
  wire NMP_PrepareWriteReq_and_61_enex5;
  wire NMP_PrepareWriteReq_and_62_enex5;
  wire rva_out_reg_data_and_102_enex5;
  wire rva_out_reg_data_and_103_enex5;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_3_enex5;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_1_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_enex5;
  wire NMP_ComputeRMSNormalize_for_and_145_enex5;
  wire NMP_ComputeRMSNormalize_for_and_146_enex5;
  wire NMP_ComputeRMSNormalize_for_and_147_enex5;
  wire NMP_ComputeRMSNormalize_for_and_148_enex5;
  wire NMP_ComputeRMSNormalize_for_and_149_enex5;
  wire NMP_ComputeRMSNormalize_for_and_150_enex5;
  wire NMP_ComputeRMSNormalize_for_and_151_enex5;
  wire NMP_ComputeRMSNormalize_for_and_152_enex5;
  wire NMP_ComputeRMSNormalize_for_and_153_enex5;
  wire NMP_ComputeRMSNormalize_for_and_154_enex5;
  wire NMP_ComputeRMSNormalize_for_and_155_enex5;
  wire NMP_ComputeRMSNormalize_for_and_156_enex5;
  wire NMP_ComputeRMSNormalize_for_and_157_enex5;
  wire NMP_ComputeRMSNormalize_for_and_158_enex5;
  wire NMP_ComputeRMSNormalize_for_and_159_enex5;
  wire NMP_ComputeRMSNormalize_for_and_160_enex5;
  wire sum_exp_and_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_80_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_81_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_82_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_83_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_84_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_85_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_86_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_87_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_88_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_89_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_90_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_91_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_92_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_93_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_94_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_95_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_1_enex5;
  wire sum_exp_and_1_enex5;
  wire sum_exp_and_2_enex5;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_12_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_50_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_51_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_52_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_53_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_54_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_55_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_56_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_57_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_58_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_59_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_60_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_61_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_62_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_63_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_64_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_65_enex5;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_5_enex5;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_6_enex5;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_5_enex5;
  wire and_1085_enex5;
  wire NMP_RunFSM_switch_lp_and_126_enex5;
  wire NMP_ComputeSoftmaxMax_for_and_enex5;
  wire max_value_and_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_66_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_67_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_68_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_69_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_70_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_21_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_71_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_72_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_73_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_74_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_75_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_76_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_77_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_78_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_79_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_80_enex5;
  wire sum_exp_and_3_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_96_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_97_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_98_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_99_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_100_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_101_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_102_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_103_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_104_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_105_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_106_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_107_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_108_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_109_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_110_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_111_enex5;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_2_enex5;
  wire NMP_ComputeRMSNormalize_for_and_161_enex5;
  wire NMP_ComputeRMSNormalize_for_and_162_enex5;
  wire NMP_ComputeRMSNormalize_for_and_163_enex5;
  wire NMP_ComputeRMSNormalize_for_and_164_enex5;
  wire NMP_ComputeRMSNormalize_for_and_165_enex5;
  wire NMP_ComputeRMSNormalize_for_and_166_enex5;
  wire NMP_ComputeRMSNormalize_for_and_167_enex5;
  wire NMP_ComputeRMSNormalize_for_and_168_enex5;
  wire NMP_ComputeRMSNormalize_for_and_169_enex5;
  wire NMP_ComputeRMSNormalize_for_and_170_enex5;
  wire NMP_ComputeRMSNormalize_for_and_171_enex5;
  wire NMP_ComputeRMSNormalize_for_and_172_enex5;
  wire NMP_ComputeRMSNormalize_for_and_173_enex5;
  wire NMP_ComputeRMSNormalize_for_and_174_enex5;
  wire NMP_ComputeRMSNormalize_for_and_175_enex5;
  wire NMP_ComputeRMSNormalize_for_and_176_enex5;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_4_enex5;
  wire rva_out_reg_data_and_104_enex5;
  wire rva_out_reg_data_and_105_enex5;
  wire sum_exp_and_4_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_8_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_9_enex5;
  wire max_value_and_9_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_112_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_113_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_114_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_115_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_116_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_117_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_118_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_119_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_120_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_121_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_122_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_123_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_124_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_125_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_126_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_127_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_81_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_82_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_83_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_84_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_85_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_86_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_87_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_88_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_89_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_90_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_91_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_92_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_93_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_94_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_95_enex5;
  wire NMP_ComputeRMSNormalize_for_and_177_enex5;
  wire NMP_ComputeRMSNormalize_for_and_178_enex5;
  wire NMP_ComputeRMSNormalize_for_and_179_enex5;
  wire NMP_ComputeRMSNormalize_for_and_180_enex5;
  wire NMP_ComputeRMSNormalize_for_and_181_enex5;
  wire NMP_ComputeRMSNormalize_for_and_182_enex5;
  wire NMP_ComputeRMSNormalize_for_and_183_enex5;
  wire NMP_ComputeRMSNormalize_for_and_184_enex5;
  wire NMP_ComputeRMSNormalize_for_and_185_enex5;
  wire NMP_ComputeRMSNormalize_for_and_186_enex5;
  wire NMP_ComputeRMSNormalize_for_and_187_enex5;
  wire NMP_ComputeRMSNormalize_for_and_188_enex5;
  wire NMP_ComputeRMSNormalize_for_and_189_enex5;
  wire NMP_ComputeRMSNormalize_for_and_190_enex5;
  wire NMP_ComputeRMSNormalize_for_and_191_enex5;
  wire NMP_ComputeRMSNormalize_for_and_192_enex5;
  wire NMP_PrepareReadReq_and_56_enex5;
  wire rva_out_reg_data_and_106_enex5;
  wire rva_out_reg_data_and_107_enex5;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_13_enex5;
  wire operator_40_0_false_AC_TRN_AC_WRAP_1_and_enex5;
  wire sum_exp_and_5_enex5;
  wire NMP_RunFSM_switch_lp_and_342_enex5;
  wire NMP_PrepareWriteReq_and_63_enex5;
  wire NMP_PrepareWriteReq_and_64_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_128_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_129_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_130_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_131_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_132_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_133_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_134_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_135_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_136_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_137_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_138_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_139_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_140_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_141_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_142_enex5;
  wire NMP_ComputeSoftmaxNormalize_for_and_143_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_96_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_97_enex5;
  wire NMP_ComputeSoftmaxExp_for_and_98_enex5;
  wire NMP_ComputeRMSNormalize_for_and_193_enex5;
  wire NMP_ComputeRMSNormalize_for_and_194_enex5;
  wire NMP_ComputeRMSNormalize_for_and_195_enex5;
  wire NMP_ComputeRMSNormalize_for_and_196_enex5;
  wire NMP_ComputeRMSNormalize_for_and_197_enex5;
  wire NMP_ComputeRMSNormalize_for_and_198_enex5;
  wire NMP_ComputeRMSNormalize_for_and_199_enex5;
  wire NMP_ComputeRMSNormalize_for_and_200_enex5;
  wire NMP_ComputeRMSNormalize_for_and_201_enex5;
  wire NMP_ComputeRMSNormalize_for_and_202_enex5;
  wire NMP_ComputeRMSNormalize_for_and_203_enex5;
  wire NMP_ComputeRMSNormalize_for_and_204_enex5;
  wire NMP_ComputeRMSNormalize_for_and_205_enex5;
  wire NMP_ComputeRMSNormalize_for_and_206_enex5;
  wire NMP_ComputeRMSNormalize_for_and_207_enex5;
  wire NMP_ComputeRMSNormalize_for_and_208_enex5;
  wire NMP_PrepareReadReq_and_57_enex5;
  wire rva_out_reg_data_and_108_enex5;
  wire rva_out_reg_data_and_109_enex5;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_14_enex5;
  wire max_value_and_10_enex5;
  wire NMP_ComputeRMSNormalize_for_and_209_enex5;
  wire NMP_ComputeRMSNormalize_for_and_210_enex5;
  wire NMP_ComputeRMSNormalize_for_and_211_enex5;
  wire NMP_ComputeRMSNormalize_for_and_212_enex5;
  wire NMP_ComputeRMSNormalize_for_and_213_enex5;
  wire NMP_ComputeRMSNormalize_for_and_214_enex5;
  wire NMP_ComputeRMSNormalize_for_and_215_enex5;
  wire NMP_ComputeRMSNormalize_for_and_216_enex5;
  wire NMP_ComputeRMSNormalize_for_and_217_enex5;
  wire NMP_ComputeRMSNormalize_for_and_218_enex5;
  wire NMP_ComputeRMSNormalize_for_and_219_enex5;
  wire NMP_ComputeRMSNormalize_for_and_220_enex5;
  wire NMP_ComputeRMSNormalize_for_and_221_enex5;
  wire NMP_ComputeRMSNormalize_for_and_222_enex5;
  wire NMP_ComputeRMSNormalize_for_and_223_enex5;
  wire NMP_ComputeRMSNormalize_for_and_224_enex5;
  wire rva_out_reg_data_and_110_enex5;
  wire rva_out_reg_data_and_111_enex5;
  wire NMP_ComputeRMSNormalize_for_and_225_enex5;
  wire NMP_ComputeRMSNormalize_for_and_226_enex5;
  wire NMP_ComputeRMSNormalize_for_and_227_enex5;
  wire NMP_ComputeRMSNormalize_for_and_228_enex5;
  wire NMP_ComputeRMSNormalize_for_and_229_enex5;
  wire NMP_ComputeRMSNormalize_for_and_230_enex5;
  wire NMP_ComputeRMSNormalize_for_and_231_enex5;
  wire NMP_ComputeRMSNormalize_for_and_232_enex5;
  wire NMP_ComputeRMSNormalize_for_and_233_enex5;
  wire NMP_ComputeRMSNormalize_for_and_234_enex5;
  wire NMP_ComputeRMSNormalize_for_and_235_enex5;
  wire NMP_ComputeRMSNormalize_for_and_236_enex5;
  wire NMP_ComputeRMSNormalize_for_and_237_enex5;
  wire NMP_ComputeRMSNormalize_for_and_238_enex5;
  wire NMP_ComputeRMSNormalize_for_and_239_enex5;
  wire NMP_ComputeRMSNormalize_for_and_240_enex5;
  wire rva_out_reg_data_and_112_enex5;
  wire rva_out_reg_data_and_113_enex5;
  wire NMP_PrepareWriteReq_and_65_enex5;
  wire NMP_PrepareWriteReq_and_66_enex5;
  wire NMP_PrepareWriteReq_and_67_enex5;
  wire NMP_ComputeRMSNormalize_for_and_241_enex5;
  wire NMP_ComputeRMSNormalize_for_and_242_enex5;
  wire NMP_ComputeRMSNormalize_for_and_243_enex5;
  wire NMP_ComputeRMSNormalize_for_and_244_enex5;
  wire NMP_ComputeRMSNormalize_for_and_245_enex5;
  wire NMP_ComputeRMSNormalize_for_and_246_enex5;
  wire NMP_ComputeRMSNormalize_for_and_247_enex5;
  wire NMP_ComputeRMSNormalize_for_and_248_enex5;
  wire NMP_ComputeRMSNormalize_for_and_249_enex5;
  wire NMP_ComputeRMSNormalize_for_and_250_enex5;
  wire NMP_ComputeRMSNormalize_for_and_251_enex5;
  wire NMP_ComputeRMSNormalize_for_and_252_enex5;
  wire NMP_ComputeRMSNormalize_for_and_253_enex5;
  wire NMP_ComputeRMSNormalize_for_and_254_enex5;
  wire NMP_ComputeRMSNormalize_for_and_255_enex5;
  wire NMP_ComputeRMSNormalize_for_and_256_enex5;
  wire NMP_PrepareReadReq_and_58_enex5;
  wire NMP_PrepareReadReq_and_59_enex5;
  wire rva_out_reg_data_and_114_enex5;
  wire rva_out_reg_data_and_115_enex5;
  wire NMP_ComputeRMSNormalize_for_and_257_enex5;
  wire NMP_ComputeRMSNormalize_for_and_258_enex5;
  wire NMP_ComputeRMSNormalize_for_and_259_enex5;
  wire NMP_ComputeRMSNormalize_for_and_260_enex5;
  wire NMP_ComputeRMSNormalize_for_and_261_enex5;
  wire NMP_ComputeRMSNormalize_for_and_262_enex5;
  wire NMP_ComputeRMSNormalize_for_and_263_enex5;
  wire NMP_ComputeRMSNormalize_for_and_264_enex5;
  wire NMP_ComputeRMSNormalize_for_and_265_enex5;
  wire NMP_ComputeRMSNormalize_for_and_266_enex5;
  wire NMP_ComputeRMSNormalize_for_and_267_enex5;
  wire NMP_ComputeRMSNormalize_for_and_268_enex5;
  wire NMP_ComputeRMSNormalize_for_and_269_enex5;
  wire NMP_ComputeRMSNormalize_for_and_270_enex5;
  wire NMP_ComputeRMSNormalize_for_and_271_enex5;
  wire rva_out_reg_data_and_116_enex5;
  wire rva_out_reg_data_and_117_enex5;
  wire NMP_ComputeRMSNormalize_for_and_272_enex5;
  wire NMP_ComputeRMSNormalize_for_and_273_enex5;
  wire rva_out_reg_data_and_118_enex5;
  wire rva_out_reg_data_and_119_enex5;
  wire rva_out_reg_data_and_120_enex5;
  wire rva_out_reg_data_and_121_enex5;
  wire NMP_PrepareWriteReq_and_68_enex5;
  wire rva_out_reg_data_and_122_enex5;
  wire rva_out_reg_data_and_123_enex5;
  wire NMP_PrepareWriteReq_and_69_enex5;
  wire rva_out_reg_data_and_124_enex5;
  wire rva_out_reg_data_and_125_enex5;
  wire NMP_PrepareWriteReq_and_70_enex5;
  wire NMP_PrepareWriteReq_and_71_enex5;
  wire NMP_PrepareReadReq_and_60_enex5;
  wire rva_out_reg_data_and_126_enex5;
  wire rva_out_reg_data_and_127_enex5;
  wire NMP_PrepareWriteReq_and_72_enex5;
  wire NMP_PrepareWriteReq_and_73_enex5;
  wire NMP_PrepareReadReq_and_61_enex5;
  wire NMP_PrepareReadReq_and_62_enex5;
  wire rva_out_reg_data_and_128_enex5;
  wire rva_out_reg_data_and_129_enex5;
  wire NMP_PrepareWriteReq_and_74_enex5;
  wire NMP_PrepareWriteReq_and_75_enex5;
  wire rva_out_reg_data_and_130_enex5;
  wire rva_out_reg_data_and_131_enex5;
  wire NMP_PrepareWriteReq_and_76_enex5;
  wire NMP_PrepareWriteReq_and_77_enex5;
  wire rva_out_reg_data_and_132_enex5;
  wire rva_out_reg_data_and_133_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_3_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_4_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_5_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5;
  wire NMP_PrepareReadReq_and_63_enex5;
  wire NMP_ComputeRMSSqrtRecip_variance_and_enex5;
  wire NMP_ComputeRMSSqrtRecip_variance_and_2_enex5;
  wire NMP_PrepareReadReq_and_64_enex5;
  wire NMP_PrepareReadReq_and_65_enex5;
  wire NMP_PrepareWriteReq_and_78_enex5;
  wire NMP_PrepareWriteReq_and_79_enex5;
  wire NMP_PrepareReadReq_and_66_enex5;
  wire NMP_PrepareWriteReq_and_80_enex5;
  wire NMP_PrepareWriteReq_and_81_enex5;
  wire NMP_PrepareReadReq_and_67_enex5;
  wire NMP_PrepareWriteReq_and_82_enex5;
  wire NMP_PrepareReadReq_and_68_enex5;
  wire NMP_PrepareWriteReq_and_83_enex5;
  wire NMP_PrepareReadReq_and_69_enex5;
  wire NMP_PrepareReadReq_and_70_enex5;
  wire NMP_PrepareReadReq_and_71_enex5;
  wire NMP_PrepareReadReq_and_72_enex5;
  wire NMP_PrepareReadReq_and_73_enex5;
  wire NMP_PrepareReadReq_and_74_enex5;
  wire NMP_PrepareWriteReq_and_84_enex5;
  wire NMP_PrepareWriteReq_and_85_enex5;
  wire NMP_PrepareWriteReq_and_86_enex5;
  wire NMP_PrepareReadReq_and_75_enex5;
  wire NMP_PrepareReadReq_and_76_enex5;
  wire NMP_PrepareWriteReq_and_87_enex5;
  wire NMP_PrepareWriteReq_and_88_enex5;
  wire NMP_PrepareReadReq_and_77_enex5;
  wire NMP_PrepareWriteReq_and_89_enex5;
  wire NMP_PrepareReadReq_and_78_enex5;
  wire NMP_PrepareReadReq_and_79_enex5;
  wire NMP_PrepareWriteReq_and_90_enex5;
  wire NMP_PrepareReadReq_and_80_enex5;
  wire NMP_PrepareReadReq_and_81_enex5;
  wire NMP_PrepareWriteReq_and_91_enex5;
  wire NMP_PrepareWriteReq_and_92_enex5;
  wire NMP_PrepareWriteReq_and_93_enex5;
  wire NMP_PrepareReadReq_and_82_enex5;
  wire NMP_PrepareReadReq_and_83_enex5;
  wire NMP_PrepareWriteReq_and_94_enex5;
  wire NMP_PrepareWriteReq_and_95_enex5;
  wire NMP_PrepareReadReq_and_84_enex5;
  wire NMP_PrepareWriteReq_and_96_enex5;
  wire NMP_PrepareReadReq_and_85_enex5;
  wire NMP_PrepareWriteReq_and_97_enex5;
  wire NMP_PrepareReadReq_and_86_enex5;
  wire NMP_PrepareWriteReq_and_98_enex5;
  wire NMP_PrepareReadReq_and_87_enex5;
  wire NMP_PrepareReadReq_and_88_enex5;
  wire NMP_PrepareWriteReq_and_99_enex5;
  wire out_float_round_32_if_m_1_and_15_tmp;
  wire out_float_round_32_if_m_1_and_31_tmp;
  wire out_float_round_32_1_if_m_1_and_31_tmp;
  wire out_float_round_32_1_if_m_1_and_15_tmp;
  wire out_float_round_32_if_m_1_and_14_tmp;
  wire out_float_round_32_if_m_1_and_30_tmp;
  wire out_float_round_32_1_if_m_1_and_14_tmp;
  wire out_float_round_32_1_if_m_1_and_30_tmp;
  wire out_float_round_32_if_m_1_and_29_tmp;
  wire out_float_round_32_if_m_1_and_13_tmp;
  wire out_float_round_32_1_if_m_1_and_29_tmp;
  wire out_float_round_32_1_if_m_1_and_13_tmp;
  wire out_float_round_32_if_m_1_and_12_tmp;
  wire out_float_round_32_if_m_1_and_28_tmp;
  wire out_float_round_32_1_if_m_1_and_12_tmp;
  wire out_float_round_32_1_if_m_1_and_28_tmp;
  wire out_float_round_32_if_m_1_and_27_tmp;
  wire out_float_round_32_if_m_1_and_11_tmp;
  wire out_float_round_32_1_if_m_1_and_27_tmp;
  wire out_float_round_32_1_if_m_1_and_11_tmp;
  wire out_float_round_32_if_m_1_and_26_tmp;
  wire out_float_round_32_if_m_1_and_10_tmp;
  wire out_float_round_32_1_if_m_1_and_10_tmp;
  wire out_float_round_32_1_if_m_1_and_26_tmp;
  wire out_float_round_32_if_m_1_and_25_tmp;
  wire out_float_round_32_if_m_1_and_9_tmp;
  wire out_float_round_32_1_if_m_1_and_25_tmp;
  wire out_float_round_32_1_if_m_1_and_9_tmp;
  wire out_float_round_32_if_m_1_and_24_tmp;
  wire out_float_round_32_if_m_1_and_8_tmp;
  wire out_float_round_32_1_if_m_1_and_8_tmp;
  wire out_float_round_32_1_if_m_1_and_24_tmp;
  wire out_float_round_32_if_m_1_and_7_tmp;
  wire out_float_round_32_if_m_1_and_23_tmp;
  wire out_float_round_32_1_if_m_1_and_23_tmp;
  wire out_float_round_32_1_if_m_1_and_7_tmp;
  wire out_float_round_32_if_m_1_and_22_tmp;
  wire out_float_round_32_if_m_1_and_6_tmp;
  wire out_float_round_32_1_if_m_1_and_22_tmp;
  wire out_float_round_32_1_if_m_1_and_6_tmp;
  wire out_float_round_32_if_m_1_and_21_tmp;
  wire out_float_round_32_if_m_1_and_5_tmp;
  wire out_float_round_32_1_if_m_1_and_21_tmp;
  wire out_float_round_32_1_if_m_1_and_5_tmp;
  wire out_float_round_32_if_m_1_and_20_tmp;
  wire out_float_round_32_if_m_1_and_4_tmp;
  wire out_float_round_32_1_if_m_1_and_4_tmp;
  wire out_float_round_32_1_if_m_1_and_20_tmp;
  wire out_float_round_32_if_m_1_and_19_tmp;
  wire out_float_round_32_if_m_1_and_3_tmp;
  wire out_float_round_32_1_if_m_1_and_19_tmp;
  wire out_float_round_32_1_if_m_1_and_3_tmp;
  wire out_float_round_32_if_m_1_and_2_tmp;
  wire out_float_round_32_if_m_1_and_18_tmp;
  wire out_float_round_32_1_if_m_1_and_18_tmp;
  wire out_float_round_32_1_if_m_1_and_2_tmp;
  wire out_float_round_32_if_m_1_and_1_tmp;
  wire out_float_round_32_if_m_1_and_17_tmp;
  wire out_float_round_32_1_if_m_1_and_1_tmp;
  wire out_float_round_32_1_if_m_1_and_17_tmp;
  wire out_float_round_32_if_m_1_and_tmp;
  wire out_float_round_32_if_m_1_and_16_tmp;
  wire out_float_round_32_1_if_m_1_and_16_tmp;
  wire out_float_round_32_1_if_m_1_and_tmp;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp;
  wire NMP_ComputeSoftmaxMax_for_if_and_tmp;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_tmp;
  wire and_1082_tmp;
  wire and_1063_tmp;
  wire and_1236_itm;
  wire mux_149_itm;
  wire NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_54_itm;
  wire [25:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_52_itm;
  wire or_924_itm;
  wire max_value_mux_1_itm;
  wire [25:0] max_value_mux_2_itm;
  wire operator_8_false_acc_1_itm_9_1;
  wire operator_16_false_acc_2_itm_17;
  wire [24:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_itm_35_11_1;
  wire mux_219_cse;
  wire mux_146_cse;

  wire mux_16_nl;
  wire nor_201_nl;
  wire or_504_nl;
  wire mux_18_nl;
  wire nor_202_nl;
  wire or_508_nl;
  wire mux_19_nl;
  wire nor_203_nl;
  wire or_514_nl;
  wire mux_21_nl;
  wire nor_204_nl;
  wire or_518_nl;
  wire or_538_nl;
  wire mux_48_nl;
  wire mux_47_nl;
  wire mux_46_nl;
  wire mux_45_nl;
  wire mux_41_nl;
  wire mux_38_nl;
  wire or_536_nl;
  wire or_535_nl;
  wire mux_37_nl;
  wire mux_36_nl;
  wire mux_35_nl;
  wire mux_34_nl;
  wire mux_24_nl;
  wire mux_33_nl;
  wire mux_32_nl;
  wire mux_30_nl;
  wire nor_5_nl;
  wire mux_29_nl;
  wire mux_28_nl;
  wire or_532_nl;
  wire or_524_nl;
  wire mux_50_nl;
  wire nor_205_nl;
  wire and_893_nl;
  wire mux_79_nl;
  wire or_555_nl;
  wire mux_80_nl;
  wire or_557_nl;
  wire[39:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_33_nl;
  wire[39:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux_nl;
  wire NMP_RunFSM_switch_lp_and_7_nl;
  wire NMP_RunFSM_switch_lp_not_63_nl;
  wire rms_reciprocal_and_nl;
  wire[39:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_32_nl;
  wire[39:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux_1_nl;
  wire NMP_RunFSM_switch_lp_and_5_nl;
  wire NMP_RunFSM_switch_lp_not_49_nl;
  wire sum_exp_reciprocal_and_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_16_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_15_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_16_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_16_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_127_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_16_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_15_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_16_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_127_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_17_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_14_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_15_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_15_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_126_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_17_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_14_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_15_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_126_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_18_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_13_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_14_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_14_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_125_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_18_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_13_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_14_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_125_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_19_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_12_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_13_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_13_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_124_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_19_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_12_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_13_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_124_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_20_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_11_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_12_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_12_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_123_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_20_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_11_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_12_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_123_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_21_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_10_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_11_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_11_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_122_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_21_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_10_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_11_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_122_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_22_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_9_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_10_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_10_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_121_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_22_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_9_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_10_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_121_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_23_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_8_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_9_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_9_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_120_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_23_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_8_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_9_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_120_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_24_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_7_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_8_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_8_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_119_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_24_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_7_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_8_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_119_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_25_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_6_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_7_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_7_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_118_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_25_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_6_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_7_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_118_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_26_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_5_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_6_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_6_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_117_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_26_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_5_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_6_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_117_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_27_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_4_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_5_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_5_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_116_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_27_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_4_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_5_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_116_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_28_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_3_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_4_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_4_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_115_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_28_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_3_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_4_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_115_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_29_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_2_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_3_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_3_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_114_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_29_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_2_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_3_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_114_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_30_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_1_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_2_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_2_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_113_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_30_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_1_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_2_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_113_nl;
  wire[3:0] out_adp_set_value_ac_float_nor_31_nl;
  wire[3:0] out_adp_set_value_ac_float_else_1_else_mux_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_for_1_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_for_1_out_adp_set_value_ac_float_else_1_else_if_acc_nl;
  wire operator_5_true_not_112_nl;
  wire[3:0] out_adp_set_value_ac_float_1_nor_31_nl;
  wire[3:0] out_adp_set_value_ac_float_1_else_1_else_mux_nl;
  wire[3:0] NMP_ConvertOutputToAdpfloat_1_for_1_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire[4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl;
  wire operator_5_true_1_not_112_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_30_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_29_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_29_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_27_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_28_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_27_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_23_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_26_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_21_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_25_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_19_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_24_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_17_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_23_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_15_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_22_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_21_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_11_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_20_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_9_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_19_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_7_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_18_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_5_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_17_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_3_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_16_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_31_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_30_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_29_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_29_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_27_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_28_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_25_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_27_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_23_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_26_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_21_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_25_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_19_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_24_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_17_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_23_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_15_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_22_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_13_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_21_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_11_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_20_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_9_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_19_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_7_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_18_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_5_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_17_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_3_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_16_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl;
  wire[4:0] out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_1_nl;
  wire[4:0] NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[5:0] nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_51_nl;
  wire NMP_RunFSM_switch_lp_not_64_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_50_nl;
  wire NMP_RunFSM_switch_lp_not_65_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_49_nl;
  wire NMP_RunFSM_switch_lp_not_66_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_48_nl;
  wire NMP_RunFSM_switch_lp_not_67_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_47_nl;
  wire NMP_RunFSM_switch_lp_not_68_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_46_nl;
  wire NMP_RunFSM_switch_lp_not_69_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_45_nl;
  wire NMP_RunFSM_switch_lp_not_70_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_44_nl;
  wire NMP_RunFSM_switch_lp_not_71_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_43_nl;
  wire NMP_RunFSM_switch_lp_not_72_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_42_nl;
  wire NMP_RunFSM_switch_lp_not_73_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_41_nl;
  wire NMP_RunFSM_switch_lp_not_74_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_40_nl;
  wire NMP_RunFSM_switch_lp_not_75_nl;
  wire[26:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_39_nl;
  wire NMP_RunFSM_switch_lp_not_76_nl;
  wire NMP_RunFSM_switch_lp_mux_32_nl;
  wire mux_277_nl;
  wire NMP_RunFSM_switch_lp_or_41_nl;
  wire NMP_RunFSM_switch_lp_not_77_nl;
  wire NMP_RunFSM_switch_lp_not_78_nl;
  wire NMP_RunFSM_switch_lp_not_51_nl;
  wire[15:0] operator_16_false_acc_2_nl;
  wire[16:0] nl_operator_16_false_acc_2_nl;
  wire mux_222_nl;
  wire mux_101_nl;
  wire mux_129_nl;
  wire or_813_nl;
  wire mux_212_nl;
  wire mux_211_nl;
  wire or_877_nl;
  wire or_875_nl;
  wire mux_210_nl;
  wire mux_209_nl;
  wire mux_208_nl;
  wire mux_207_nl;
  wire mux_206_nl;
  wire mux_205_nl;
  wire mux_204_nl;
  wire mux_203_nl;
  wire mux_202_nl;
  wire mux_201_nl;
  wire and_896_nl;
  wire and_897_nl;
  wire mux_199_nl;
  wire and_673_nl;
  wire mux_197_nl;
  wire nor_211_nl;
  wire mux_196_nl;
  wire nand_18_nl;
  wire mux_195_nl;
  wire mux_193_nl;
  wire mux_192_nl;
  wire mux_191_nl;
  wire nor_212_nl;
  wire mux_186_nl;
  wire nor_213_nl;
  wire mux_184_nl;
  wire or_850_nl;
  wire and_901_nl;
  wire mux_181_nl;
  wire and_902_nl;
  wire mux_180_nl;
  wire mux_179_nl;
  wire and_903_nl;
  wire and_904_nl;
  wire mux_138_nl;
  wire mux_137_nl;
  wire mux_136_nl;
  wire mux_135_nl;
  wire mux_134_nl;
  wire mux_133_nl;
  wire mux_132_nl;
  wire mux_128_nl;
  wire mux_127_nl;
  wire mux_126_nl;
  wire mux_124_nl;
  wire mux_123_nl;
  wire mux_278_nl;
  wire mux_122_nl;
  wire or_811_nl;
  wire mux_121_nl;
  wire or_809_nl;
  wire mux_120_nl;
  wire mux_119_nl;
  wire mux_118_nl;
  wire mux_117_nl;
  wire mux_116_nl;
  wire mux_115_nl;
  wire mux_113_nl;
  wire mux_112_nl;
  wire mux_103_nl;
  wire or_790_nl;
  wire mux_82_nl;
  wire mux_81_nl;
  wire or_784_nl;
  wire and_889_nl;
  wire mux_281_nl;
  wire and_671_nl;
  wire mux_178_nl;
  wire mux_177_nl;
  wire mux_176_nl;
  wire mux_175_nl;
  wire mux_174_nl;
  wire mux_173_nl;
  wire mux_172_nl;
  wire mux_171_nl;
  wire mux_170_nl;
  wire mux_169_nl;
  wire mux_168_nl;
  wire mux_167_nl;
  wire mux_166_nl;
  wire mux_164_nl;
  wire mux_163_nl;
  wire mux_162_nl;
  wire or_836_nl;
  wire mux_160_nl;
  wire mux_159_nl;
  wire mux_158_nl;
  wire mux_157_nl;
  wire mux_155_nl;
  wire mux_154_nl;
  wire mux_153_nl;
  wire mux_282_nl;
  wire and_894_nl;
  wire or_830_nl;
  wire or_820_nl;
  wire mux_141_nl;
  wire nand_2_nl;
  wire or_815_nl;
  wire[39:0] NMP_ComputeRMSSumSq_for_acc_nl;
  wire[43:0] nl_NMP_ComputeRMSSumSq_for_acc_nl;
  wire[39:0] NMP_ComputeRMSSumSq_for_acc_3_nl;
  wire[42:0] nl_NMP_ComputeRMSSumSq_for_acc_3_nl;
  wire NMP_PrepareReadReq_or_nl;
  wire mux_15_nl;
  wire nor_66_nl;
  wire nor_67_nl;
  wire nmp_config_ConfigRead_not_12_nl;
  wire nmp_config_ConfigRead_not_10_nl;
  wire nmp_config_ConfigRead_not_9_nl;
  wire nmp_config_ConfigRead_not_6_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_45_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_45_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_32_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_32_nl;
  wire operator_5_true_not_110_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_32_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_32_nl;
  wire operator_5_true_1_not_110_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_15_nl;
  wire out_adp_set_value_ac_float_mux_75_nl;
  wire operator_5_true_mux_31_nl;
  wire or_668_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_15_nl;
  wire out_adp_set_value_ac_float_1_mux_75_nl;
  wire operator_5_true_1_mux_31_nl;
  wire or_766_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_33_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_33_nl;
  wire operator_5_true_not_80_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_33_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_33_nl;
  wire operator_5_true_1_not_80_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_nl;
  wire out_adp_set_value_ac_float_mux_nl;
  wire operator_5_true_mux_1_nl;
  wire or_578_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_nl;
  wire out_adp_set_value_ac_float_1_mux_nl;
  wire operator_5_true_1_mux_1_nl;
  wire or_676_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_42_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_42_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_34_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_34_nl;
  wire operator_5_true_not_108_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_34_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_34_nl;
  wire operator_5_true_1_not_108_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_14_nl;
  wire out_adp_set_value_ac_float_mux_70_nl;
  wire operator_5_true_mux_29_nl;
  wire or_662_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_14_nl;
  wire out_adp_set_value_ac_float_1_mux_70_nl;
  wire operator_5_true_1_mux_29_nl;
  wire or_760_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_35_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_35_nl;
  wire operator_5_true_not_82_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_35_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_35_nl;
  wire operator_5_true_1_not_82_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_1_nl;
  wire out_adp_set_value_ac_float_mux_5_nl;
  wire operator_5_true_mux_3_nl;
  wire or_584_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_1_nl;
  wire out_adp_set_value_ac_float_1_mux_5_nl;
  wire operator_5_true_1_mux_3_nl;
  wire or_682_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_3_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_3_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_39_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_39_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_36_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_36_nl;
  wire operator_5_true_not_106_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_36_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_36_nl;
  wire operator_5_true_1_not_106_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_13_nl;
  wire out_adp_set_value_ac_float_mux_65_nl;
  wire operator_5_true_mux_27_nl;
  wire or_656_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_13_nl;
  wire out_adp_set_value_ac_float_1_mux_65_nl;
  wire operator_5_true_1_mux_27_nl;
  wire or_754_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_37_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_37_nl;
  wire operator_5_true_not_84_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_37_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_37_nl;
  wire operator_5_true_1_not_84_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_2_nl;
  wire out_adp_set_value_ac_float_mux_10_nl;
  wire operator_5_true_mux_5_nl;
  wire or_590_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_2_nl;
  wire out_adp_set_value_ac_float_1_mux_10_nl;
  wire operator_5_true_1_mux_5_nl;
  wire or_688_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_6_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_6_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_36_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_36_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_38_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_38_nl;
  wire operator_5_true_not_104_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_38_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_38_nl;
  wire operator_5_true_1_not_104_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_12_nl;
  wire out_adp_set_value_ac_float_mux_60_nl;
  wire operator_5_true_mux_25_nl;
  wire or_650_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_12_nl;
  wire out_adp_set_value_ac_float_1_mux_60_nl;
  wire operator_5_true_1_mux_25_nl;
  wire or_748_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_39_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_39_nl;
  wire operator_5_true_not_86_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_39_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_39_nl;
  wire operator_5_true_1_not_86_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_3_nl;
  wire out_adp_set_value_ac_float_mux_15_nl;
  wire operator_5_true_mux_7_nl;
  wire or_596_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_3_nl;
  wire out_adp_set_value_ac_float_1_mux_15_nl;
  wire operator_5_true_1_mux_7_nl;
  wire or_694_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_9_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_9_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_33_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_33_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_40_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_40_nl;
  wire operator_5_true_not_102_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_40_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_40_nl;
  wire operator_5_true_1_not_102_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_11_nl;
  wire out_adp_set_value_ac_float_mux_55_nl;
  wire operator_5_true_mux_23_nl;
  wire or_644_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_11_nl;
  wire out_adp_set_value_ac_float_1_mux_55_nl;
  wire operator_5_true_1_mux_23_nl;
  wire or_742_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_41_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_41_nl;
  wire operator_5_true_not_88_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_41_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_41_nl;
  wire operator_5_true_1_not_88_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_4_nl;
  wire out_adp_set_value_ac_float_mux_20_nl;
  wire operator_5_true_mux_9_nl;
  wire or_602_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_4_nl;
  wire out_adp_set_value_ac_float_1_mux_20_nl;
  wire operator_5_true_1_mux_9_nl;
  wire or_700_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_12_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_12_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_30_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_30_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_42_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_42_nl;
  wire operator_5_true_not_100_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_42_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_42_nl;
  wire operator_5_true_1_not_100_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_10_nl;
  wire out_adp_set_value_ac_float_mux_50_nl;
  wire operator_5_true_mux_21_nl;
  wire or_638_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_10_nl;
  wire out_adp_set_value_ac_float_1_mux_50_nl;
  wire operator_5_true_1_mux_21_nl;
  wire or_736_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_43_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_43_nl;
  wire operator_5_true_not_90_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_43_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_43_nl;
  wire operator_5_true_1_not_90_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_5_nl;
  wire out_adp_set_value_ac_float_mux_25_nl;
  wire operator_5_true_mux_11_nl;
  wire or_608_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_5_nl;
  wire out_adp_set_value_ac_float_1_mux_25_nl;
  wire operator_5_true_1_mux_11_nl;
  wire or_706_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_15_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_15_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_27_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_27_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_44_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_44_nl;
  wire operator_5_true_not_98_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_44_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_44_nl;
  wire operator_5_true_1_not_98_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_9_nl;
  wire out_adp_set_value_ac_float_mux_45_nl;
  wire operator_5_true_mux_19_nl;
  wire or_632_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_9_nl;
  wire out_adp_set_value_ac_float_1_mux_45_nl;
  wire operator_5_true_1_mux_19_nl;
  wire or_730_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_45_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_45_nl;
  wire operator_5_true_not_92_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_45_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_45_nl;
  wire operator_5_true_1_not_92_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_6_nl;
  wire out_adp_set_value_ac_float_mux_30_nl;
  wire operator_5_true_mux_13_nl;
  wire or_614_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_6_nl;
  wire out_adp_set_value_ac_float_1_mux_30_nl;
  wire operator_5_true_1_mux_13_nl;
  wire or_712_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_18_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_18_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_24_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_24_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_46_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_46_nl;
  wire operator_5_true_not_96_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_46_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_46_nl;
  wire operator_5_true_1_not_96_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_8_nl;
  wire out_adp_set_value_ac_float_mux_40_nl;
  wire operator_5_true_mux_17_nl;
  wire or_626_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_8_nl;
  wire out_adp_set_value_ac_float_1_mux_40_nl;
  wire operator_5_true_1_mux_17_nl;
  wire or_724_nl;
  wire[1:0] out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_47_nl;
  wire[1:0] out_adp_set_value_ac_float_nor_47_nl;
  wire operator_5_true_not_94_nl;
  wire[1:0] out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_47_nl;
  wire[1:0] out_adp_set_value_ac_float_1_nor_47_nl;
  wire operator_5_true_1_not_94_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_7_nl;
  wire out_adp_set_value_ac_float_mux_35_nl;
  wire operator_5_true_mux_15_nl;
  wire or_620_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_7_nl;
  wire out_adp_set_value_ac_float_1_mux_35_nl;
  wire operator_5_true_1_mux_15_nl;
  wire or_718_nl;
  wire out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_21_nl;
  wire out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_21_nl;
  wire[7:0] mux_258_nl;
  wire[7:0] while_while_while_or_nl;
  wire or_922_nl;
  wire nor_266_nl;
  wire[9:0] operator_8_false_acc_1_nl;
  wire[11:0] nl_operator_8_false_acc_1_nl;
  wire NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux1h_3_nl;
  wire NMP_RunFSM_switch_lp_and_24_nl;
  wire[25:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux_2_nl;
  wire NMP_RunFSM_switch_lp_not_80_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_31_nl;
  wire NMP_RunFSM_switch_lp_not_81_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_30_nl;
  wire NMP_RunFSM_switch_lp_not_82_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_29_nl;
  wire NMP_RunFSM_switch_lp_not_83_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_28_nl;
  wire NMP_RunFSM_switch_lp_not_84_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_27_nl;
  wire NMP_RunFSM_switch_lp_not_85_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_26_nl;
  wire NMP_RunFSM_switch_lp_not_86_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_25_nl;
  wire NMP_RunFSM_switch_lp_not_87_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_24_nl;
  wire NMP_RunFSM_switch_lp_not_88_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_23_nl;
  wire NMP_RunFSM_switch_lp_not_89_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_22_nl;
  wire NMP_RunFSM_switch_lp_not_90_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_21_nl;
  wire NMP_RunFSM_switch_lp_not_91_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_20_nl;
  wire NMP_RunFSM_switch_lp_not_92_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_19_nl;
  wire NMP_RunFSM_switch_lp_not_93_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_18_nl;
  wire NMP_RunFSM_switch_lp_not_94_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_17_nl;
  wire NMP_RunFSM_switch_lp_not_95_nl;
  wire[31:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_55_nl;
  wire NMP_RunFSM_switch_lp_not_57_nl;
  wire[35:0] NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_35_nl;
  wire NMP_RunFSM_switch_lp_not_25_nl;
  wire or_927_nl;
  wire NMP_RunFSM_switch_lp_mux1h_74_nl;
  wire NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_25_nl;
  wire NMP_RunFSM_switch_lp_mux1h_72_nl;
  wire NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_24_nl;
  wire NMP_RunFSM_switch_lp_mux_51_nl;
  wire[17:0] operator_16_false_acc_2_nl_1;
  wire[19:0] nl_operator_16_false_acc_2_nl_1;
  wire[35:0] ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_nl;
  wire[36:0] nl_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_60_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_64_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_56_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_4_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_52_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_8_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_48_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_12_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_44_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_16_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_40_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_20_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_36_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_24_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_32_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_28_nl;
  wire while_mux_1001_nl;
  wire max_value_and_11_nl;
  wire nand_3_nl;
  wire nand_nl;
  wire mux_5_nl;
  wire nor_45_nl;
  wire nor_46_nl;
  wire nor_79_nl;
  wire or_509_nl;
  wire nor_80_nl;
  wire or_519_nl;
  wire mux_280_nl;
  wire or_799_nl;
  wire mux_98_nl;
  wire nor_16_nl;
  wire or_819_nl;
  wire or_818_nl;
  wire or_823_nl;
  wire or_827_nl;
  wire mux_8_nl;
  wire nand_5_nl;
  wire nor_1_nl;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_nl;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_1_nl;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_2_nl;
  wire ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_3_nl;
  wire mux_10_nl;
  wire mux_9_nl;
  wire or_452_nl;
  wire ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_nl;
  wire[1:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_8_nl;
  wire[1:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux1h_60_nl;
  wire and_833_nl;
  wire and_836_nl;
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_not_3_nl;
  wire mux_11_nl;
  wire nor_54_nl;
  wire nor_55_nl;
  wire[1:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_4_nl;
  wire[1:0] ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux1h_59_nl;
  wire ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_nand_nl;
  wire mux_12_nl;
  wire NMP_PrepareWriteReq_and_nl;
  wire NMP_PrepareWriteReq_and_1_nl;
  wire NMP_PrepareWriteReq_and_2_nl;
  wire NMP_PrepareWriteReq_and_3_nl;
  wire mux_13_nl;
  wire NMP_PrepareReadReq_and_2_nl;
  wire NMP_PrepareReadReq_and_3_nl;
  wire NMP_PrepareReadReq_and_4_nl;
  wire NMP_PrepareReadReq_and_5_nl;
  wire mux_14_nl;
  wire and_880_nl;
  wire nmp_config_ConfigRead_nmp_config_ConfigRead_and_7_nl;
  wire[1:0] nmp_config_ConfigRead_nmp_config_ConfigRead_and_12_nl;
  wire nmp_config_ConfigRead_not_13_nl;
  wire[5:0] NMP_PrepareWriteReq_NMP_PrepareWriteReq_mux1h_1_nl;
  wire NMP_PrepareWriteReq_not_6_nl;
  wire[5:0] NMP_PrepareReadReq_NMP_PrepareReadReq_mux1h_1_nl;
  wire NMP_PrepareReadReq_not_6_nl;
  wire mux_273_nl;
  wire mux_272_nl;
  wire mux_271_nl;
  wire and_1081_nl;
  wire and_1080_nl;
  wire and_1079_nl;
  wire nand_21_nl;
  wire mux_269_nl;
  wire nor_294_nl;
  wire mux_268_nl;
  wire mux_267_nl;
  wire or_976_nl;
  wire or_975_nl;
  wire mux_266_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[10:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_mux_2_nl;
  wire[9:0] ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_mux_nl;
  wire [25:0] nl_operator_40_16_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_mux_2_nl
      = MUX_v_11_2_2(ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_psp_sva,
      (ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_qif_ac_fixed_cctor_20_0_sva_1[20:10]),
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_4_39);
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_mux_nl
      = MUX_v_10_2_2(ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1_9_0,
      (ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_qif_ac_fixed_cctor_20_0_sva_1[9:0]),
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_4_39);
  assign nl_operator_40_16_true_AC_TRN_AC_WRAP_rshift_rg_a = {ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_4_39
      , ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_mux_2_nl
      , ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_mux_nl
      , 4'b0000};
  wire [24:0] nl_operator_40_16_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_operator_40_16_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_itm
      , ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TR000000
      , 4'b0000};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_75_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_15_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_77_nl;
  wire[3:0] in_adp_to_ac_float_mux_166_nl;
  wire in_adp_is_zero_aelse_not_159_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_75_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[127])
      & (~ in_adp_is_zero_land_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_15_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[127])))) |
      in_adp_is_zero_land_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_166_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[123:120]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[127]);
  assign in_adp_is_zero_aelse_not_159_nl = ~ in_adp_is_zero_land_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_77_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_166_nl,
      in_adp_is_zero_aelse_not_159_nl);
  assign nl_NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_75_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_15_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_77_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_78_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_16_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_16_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_158_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_79_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_16_operator_4_false_acc_1_nl = 4'b1011 +
      conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_16_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_16_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_158_nl = ~ in_adp_is_zero_land_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_78_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_16_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_158_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_79_nl = (in_adp_to_ac_float_acc_sdt_sva_1[0])
      & (~ in_adp_is_zero_land_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_78_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_79_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_70_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_14_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_72_nl;
  wire[3:0] in_adp_to_ac_float_mux_155_nl;
  wire in_adp_is_zero_aelse_not_156_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_70_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[119])
      & (~ in_adp_is_zero_land_15_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_14_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_15_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[119])))) |
      in_adp_is_zero_land_15_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_155_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[115:112]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_15_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[119]);
  assign in_adp_is_zero_aelse_not_156_nl = ~ in_adp_is_zero_land_15_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_72_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_155_nl,
      in_adp_is_zero_aelse_not_156_nl);
  assign nl_NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_70_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_14_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_72_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_73_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_15_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_15_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_155_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_74_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_15_operator_4_false_acc_1_nl = 4'b1011 +
      conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_15_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_15_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_15_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_155_nl = ~ in_adp_is_zero_land_15_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_73_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_15_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_155_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_74_nl = (in_adp_to_ac_float_acc_sdt_15_sva_1[0])
      & (~ in_adp_is_zero_land_15_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_73_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_74_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_65_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_13_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_67_nl;
  wire[3:0] in_adp_to_ac_float_mux_144_nl;
  wire in_adp_is_zero_aelse_not_153_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_65_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[111])
      & (~ in_adp_is_zero_land_14_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_13_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_14_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[111])))) |
      in_adp_is_zero_land_14_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_144_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[107:104]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_14_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[111]);
  assign in_adp_is_zero_aelse_not_153_nl = ~ in_adp_is_zero_land_14_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_67_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_144_nl,
      in_adp_is_zero_aelse_not_153_nl);
  assign nl_NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_65_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_13_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_67_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_68_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_14_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_14_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_152_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_69_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_14_operator_4_false_acc_1_nl = 4'b1011 +
      conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_14_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_14_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_14_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_152_nl = ~ in_adp_is_zero_land_14_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_68_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_14_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_152_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_69_nl = (in_adp_to_ac_float_acc_sdt_14_sva_1[0])
      & (~ in_adp_is_zero_land_14_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_68_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_69_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_60_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_12_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_62_nl;
  wire[3:0] in_adp_to_ac_float_mux_133_nl;
  wire in_adp_is_zero_aelse_not_150_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_60_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[103])
      & (~ in_adp_is_zero_land_13_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_12_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_13_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[103])))) |
      in_adp_is_zero_land_13_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_133_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[99:96]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_13_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[103]);
  assign in_adp_is_zero_aelse_not_150_nl = ~ in_adp_is_zero_land_13_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_62_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_133_nl,
      in_adp_is_zero_aelse_not_150_nl);
  assign nl_NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_60_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_12_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_62_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_63_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_13_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_13_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_149_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_64_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_13_operator_4_false_acc_1_nl = 4'b1011 +
      conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_13_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_13_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_13_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_149_nl = ~ in_adp_is_zero_land_13_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_63_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_13_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_149_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_64_nl = (in_adp_to_ac_float_acc_sdt_13_sva_1[0])
      & (~ in_adp_is_zero_land_13_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_63_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_64_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_55_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_11_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_57_nl;
  wire[3:0] in_adp_to_ac_float_mux_122_nl;
  wire in_adp_is_zero_aelse_not_147_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_55_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[95])
      & (~ in_adp_is_zero_land_12_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_11_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_12_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[95])))) |
      in_adp_is_zero_land_12_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_122_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[91:88]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_12_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[95]);
  assign in_adp_is_zero_aelse_not_147_nl = ~ in_adp_is_zero_land_12_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_57_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_122_nl,
      in_adp_is_zero_aelse_not_147_nl);
  assign nl_NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_55_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_11_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_57_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_58_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_12_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_12_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_146_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_59_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_12_operator_4_false_acc_1_nl = 4'b1011 +
      conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_12_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_12_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_12_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_146_nl = ~ in_adp_is_zero_land_12_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_58_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_12_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_146_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_59_nl = (in_adp_to_ac_float_acc_sdt_12_sva_1[0])
      & (~ in_adp_is_zero_land_12_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_58_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_59_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_50_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_10_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_52_nl;
  wire[3:0] in_adp_to_ac_float_mux_111_nl;
  wire in_adp_is_zero_aelse_not_144_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_50_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[87])
      & (~ in_adp_is_zero_land_11_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_10_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_11_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[87])))) |
      in_adp_is_zero_land_11_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_111_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[83:80]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_11_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[87]);
  assign in_adp_is_zero_aelse_not_144_nl = ~ in_adp_is_zero_land_11_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_52_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_111_nl,
      in_adp_is_zero_aelse_not_144_nl);
  assign nl_NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_50_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_10_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_52_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_53_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_11_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_11_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_143_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_54_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_11_operator_4_false_acc_1_nl = 4'b1011 +
      conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_11_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_11_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_11_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_143_nl = ~ in_adp_is_zero_land_11_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_53_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_11_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_143_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_54_nl = (in_adp_to_ac_float_acc_sdt_11_sva_1[0])
      & (~ in_adp_is_zero_land_11_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_53_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_54_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_45_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_9_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_47_nl;
  wire[3:0] in_adp_to_ac_float_mux_100_nl;
  wire in_adp_is_zero_aelse_not_141_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_45_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[79])
      & (~ in_adp_is_zero_land_10_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_9_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_10_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[79])))) |
      in_adp_is_zero_land_10_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_100_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[75:72]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_10_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[79]);
  assign in_adp_is_zero_aelse_not_141_nl = ~ in_adp_is_zero_land_10_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_47_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_100_nl,
      in_adp_is_zero_aelse_not_141_nl);
  assign nl_NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_45_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_9_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_47_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_48_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_10_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_10_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_140_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_49_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_10_operator_4_false_acc_1_nl = 4'b1011 +
      conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_10_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_10_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_10_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_140_nl = ~ in_adp_is_zero_land_10_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_48_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_10_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_140_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_49_nl = (in_adp_to_ac_float_acc_sdt_10_sva_1[0])
      & (~ in_adp_is_zero_land_10_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_48_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_49_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_40_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_8_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_42_nl;
  wire[3:0] in_adp_to_ac_float_mux_89_nl;
  wire in_adp_is_zero_aelse_not_138_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_40_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[71])
      & (~ in_adp_is_zero_land_9_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_8_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_9_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[71])))) |
      in_adp_is_zero_land_9_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_89_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[67:64]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_9_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[71]);
  assign in_adp_is_zero_aelse_not_138_nl = ~ in_adp_is_zero_land_9_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_42_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_89_nl,
      in_adp_is_zero_aelse_not_138_nl);
  assign nl_NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_40_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_8_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_42_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_43_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_9_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_9_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_137_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_44_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_9_operator_4_false_acc_1_nl = 4'b1011 + conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_9_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_9_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_9_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_137_nl = ~ in_adp_is_zero_land_9_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_43_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_9_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_137_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_44_nl = (in_adp_to_ac_float_acc_sdt_9_sva_1[0])
      & (~ in_adp_is_zero_land_9_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_43_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_44_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_35_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_7_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_37_nl;
  wire[3:0] in_adp_to_ac_float_mux_78_nl;
  wire in_adp_is_zero_aelse_not_135_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_35_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[63])
      & (~ in_adp_is_zero_land_8_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_7_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_8_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[63])))) |
      in_adp_is_zero_land_8_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_78_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[59:56]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_8_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[63]);
  assign in_adp_is_zero_aelse_not_135_nl = ~ in_adp_is_zero_land_8_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_37_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_78_nl,
      in_adp_is_zero_aelse_not_135_nl);
  assign nl_NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_35_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_7_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_37_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_38_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_8_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_8_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_134_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_39_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_8_operator_4_false_acc_1_nl = 4'b1011 + conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_8_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_8_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_8_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_134_nl = ~ in_adp_is_zero_land_8_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_38_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_8_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_134_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_39_nl = (in_adp_to_ac_float_acc_sdt_8_sva_1[0])
      & (~ in_adp_is_zero_land_8_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_38_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_39_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_30_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_6_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_32_nl;
  wire[3:0] in_adp_to_ac_float_mux_67_nl;
  wire in_adp_is_zero_aelse_not_132_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_30_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[55])
      & (~ in_adp_is_zero_land_7_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_6_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_7_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[55])))) |
      in_adp_is_zero_land_7_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_67_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[51:48]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_7_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[55]);
  assign in_adp_is_zero_aelse_not_132_nl = ~ in_adp_is_zero_land_7_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_32_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_67_nl,
      in_adp_is_zero_aelse_not_132_nl);
  assign nl_NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_30_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_6_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_32_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_33_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_7_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_7_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_131_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_34_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_7_operator_4_false_acc_1_nl = 4'b1011 + conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_7_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_7_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_7_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_131_nl = ~ in_adp_is_zero_land_7_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_33_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_7_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_131_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_34_nl = (in_adp_to_ac_float_acc_sdt_7_sva_1[0])
      & (~ in_adp_is_zero_land_7_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_33_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_34_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_25_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_5_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_27_nl;
  wire[3:0] in_adp_to_ac_float_mux_56_nl;
  wire in_adp_is_zero_aelse_not_129_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_25_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[47])
      & (~ in_adp_is_zero_land_6_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_5_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_6_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[47])))) |
      in_adp_is_zero_land_6_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_56_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[43:40]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_6_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[47]);
  assign in_adp_is_zero_aelse_not_129_nl = ~ in_adp_is_zero_land_6_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_27_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_56_nl,
      in_adp_is_zero_aelse_not_129_nl);
  assign nl_NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_25_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_5_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_27_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_28_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_6_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_6_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_128_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_29_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_6_operator_4_false_acc_1_nl = 4'b1011 + conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_6_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_6_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_6_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_128_nl = ~ in_adp_is_zero_land_6_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_28_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_6_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_128_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_29_nl = (in_adp_to_ac_float_acc_sdt_6_sva_1[0])
      & (~ in_adp_is_zero_land_6_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_28_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_29_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_20_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_4_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_22_nl;
  wire[3:0] in_adp_to_ac_float_mux_45_nl;
  wire in_adp_is_zero_aelse_not_126_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_20_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[39])
      & (~ in_adp_is_zero_land_5_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_4_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_5_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[39])))) |
      in_adp_is_zero_land_5_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_45_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[35:32]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_5_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[39]);
  assign in_adp_is_zero_aelse_not_126_nl = ~ in_adp_is_zero_land_5_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_22_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_45_nl,
      in_adp_is_zero_aelse_not_126_nl);
  assign nl_NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_20_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_4_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_22_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_23_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_5_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_5_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_125_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_24_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_5_operator_4_false_acc_1_nl = 4'b1011 + conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_5_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_5_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_5_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_125_nl = ~ in_adp_is_zero_land_5_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_23_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_5_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_125_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_24_nl = (in_adp_to_ac_float_acc_sdt_5_sva_1[0])
      & (~ in_adp_is_zero_land_5_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_23_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_24_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_15_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_3_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_17_nl;
  wire[3:0] in_adp_to_ac_float_mux_34_nl;
  wire in_adp_is_zero_aelse_not_123_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_15_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[31])
      & (~ in_adp_is_zero_land_4_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_3_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_4_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[31])))) |
      in_adp_is_zero_land_4_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_34_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[27:24]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_4_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[31]);
  assign in_adp_is_zero_aelse_not_123_nl = ~ in_adp_is_zero_land_4_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_17_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_34_nl,
      in_adp_is_zero_aelse_not_123_nl);
  assign nl_NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_15_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_3_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_17_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_18_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_4_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_4_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_122_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_19_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_4_operator_4_false_acc_1_nl = 4'b1011 + conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_4_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_4_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_4_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_122_nl = ~ in_adp_is_zero_land_4_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_18_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_4_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_122_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_19_nl = (in_adp_to_ac_float_acc_sdt_4_sva_1[0])
      & (~ in_adp_is_zero_land_4_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_18_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_19_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_10_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_2_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_12_nl;
  wire[3:0] in_adp_to_ac_float_mux_23_nl;
  wire in_adp_is_zero_aelse_not_120_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_10_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[23])
      & (~ in_adp_is_zero_land_3_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_2_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_3_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[23])))) |
      in_adp_is_zero_land_3_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_23_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[19:16]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_3_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[23]);
  assign in_adp_is_zero_aelse_not_120_nl = ~ in_adp_is_zero_land_3_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_12_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_23_nl,
      in_adp_is_zero_aelse_not_120_nl);
  assign nl_NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_10_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_2_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_12_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_13_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_3_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_3_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_119_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_14_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_3_operator_4_false_acc_1_nl = 4'b1011 + conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_3_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_3_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_3_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_119_nl = ~ in_adp_is_zero_land_3_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_13_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_3_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_119_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_14_nl = (in_adp_to_ac_float_acc_sdt_3_sva_1[0])
      & (~ in_adp_is_zero_land_3_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_13_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_14_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_5_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_1_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_7_nl;
  wire[3:0] in_adp_to_ac_float_mux_12_nl;
  wire in_adp_is_zero_aelse_not_117_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_5_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[15])
      & (~ in_adp_is_zero_land_2_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_1_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_2_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[15])))) |
      in_adp_is_zero_land_2_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_12_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[11:8]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_2_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[15]);
  assign in_adp_is_zero_aelse_not_117_nl = ~ in_adp_is_zero_land_2_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_7_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_12_nl,
      in_adp_is_zero_aelse_not_117_nl);
  assign nl_NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_5_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_1_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_7_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_8_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_2_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_2_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_116_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_9_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_2_operator_4_false_acc_1_nl = 4'b1011 + conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_2_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_2_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_2_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_116_nl = ~ in_adp_is_zero_land_2_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_8_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_2_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_116_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_9_nl = (in_adp_to_ac_float_acc_sdt_2_sva_1[0])
      & (~ in_adp_is_zero_land_2_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_8_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_9_nl};
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_nl;
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_2_nl;
  wire[3:0] in_adp_to_ac_float_mux_1_nl;
  wire in_adp_is_zero_aelse_not_114_nl;
  wire [21:0] nl_NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_rg_a;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_nl = (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[7])
      & (~ in_adp_is_zero_land_1_lpi_1_dfm_1);
  assign in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_nl = ~((~((in_adp_to_ac_float_if_1_ac_int_cctor_4_0_1_sva_1[4])
      | (~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[7])))) | in_adp_is_zero_land_1_lpi_1_dfm_1);
  assign in_adp_to_ac_float_mux_1_nl = MUX_v_4_2_2((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[3:0]),
      (in_adp_to_ac_float_if_1_ac_int_cctor_4_0_1_sva_1[3:0]), large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[7]);
  assign in_adp_is_zero_aelse_not_114_nl = ~ in_adp_is_zero_land_1_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_2_nl = MUX_v_4_2_2(4'b0000, in_adp_to_ac_float_mux_1_nl,
      in_adp_is_zero_aelse_not_114_nl);
  assign nl_NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_rg_a = {in_adp_to_ac_float_in_adp_to_ac_float_and_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_in_adp_to_ac_float_nor_nl , in_adp_to_ac_float_in_adp_to_ac_float_and_2_nl
      , 16'b0000000000000000};
  wire[3:0] in_adp_to_ac_float_in_adp_to_ac_float_and_3_nl;
  wire[3:0] NMP_ConvertInputToFixed_for_1_operator_4_false_acc_1_nl;
  wire[4:0] nl_NMP_ConvertInputToFixed_for_1_operator_4_false_acc_1_nl;
  wire in_adp_is_zero_aelse_not_113_nl;
  wire in_adp_to_ac_float_in_adp_to_ac_float_and_4_nl;
  wire [4:0] nl_NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_rg_s;
  assign nl_NMP_ConvertInputToFixed_for_1_operator_4_false_acc_1_nl = 4'b1011 + conv_u2s_3_4(in_adp_to_ac_float_acc_sdt_1_sva_1[3:1]);
  assign NMP_ConvertInputToFixed_for_1_operator_4_false_acc_1_nl = nl_NMP_ConvertInputToFixed_for_1_operator_4_false_acc_1_nl[3:0];
  assign in_adp_is_zero_aelse_not_113_nl = ~ in_adp_is_zero_land_1_lpi_1_dfm_1;
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_3_nl = MUX_v_4_2_2(4'b0000, NMP_ConvertInputToFixed_for_1_operator_4_false_acc_1_nl,
      in_adp_is_zero_aelse_not_113_nl);
  assign in_adp_to_ac_float_in_adp_to_ac_float_and_4_nl = (in_adp_to_ac_float_acc_sdt_1_sva_1[0])
      & (~ in_adp_is_zero_land_1_lpi_1_dfm_1);
  assign nl_NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_rg_s = {in_adp_to_ac_float_in_adp_to_ac_float_and_3_nl
      , in_adp_to_ac_float_in_adp_to_ac_float_and_4_nl};
  wire [24:0] nl_operator_40_16_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_operator_40_16_false_AC_TRN_AC_WRAP_lshift_rg_a = {ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_1_itm_1_12_9
      , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_1_itm_1_8_0
      , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_2_itm_1_10_7
      , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_2_itm_1_6_0
      , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_itm_1};
  wire[10:0] NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_16_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_62_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_63_itm_1});
  assign NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_16_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_15_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_58_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_59_itm_1});
  assign NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_15_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_14_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_54_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_55_itm_1});
  assign NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_14_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_13_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_50_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_51_itm_1});
  assign NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_13_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_12_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_46_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_47_itm_1});
  assign NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_12_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_11_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_42_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_43_itm_1});
  assign NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_11_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_10_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_38_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_39_itm_1});
  assign NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_10_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_9_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_34_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_35_itm_1});
  assign NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_9_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_8_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_30_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_31_itm_1});
  assign NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_8_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_7_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_26_itm_1
      , 1'b1 , NMP_PrepareWriteReq_asn_2_itm_7_6_0});
  assign NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_7_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_6_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_22_itm_1
      , 1'b1 , NMP_PrepareWriteReq_asn_1_itm_7_6 , NMP_PrepareWriteReq_asn_1_itm_7_5_0});
  assign NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_6_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_5_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_18_itm_1
      , 1'b1 , NMP_PrepareReadReq_asn_2_itm_7_6_0});
  assign NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_5_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_4_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_14_itm_1_2
      , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_14_itm_1_1_0
      , 1'b1 , NMP_PrepareReadReq_asn_1_itm_7_6 , NMP_PrepareReadReq_asn_1_itm_7_5_0});
  assign NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_4_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_3_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_2
      , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_1_0
      , 1'b1 , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4});
  assign NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_3_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_2_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_6_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_7_itm_1});
  assign NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_2_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001};
  wire[10:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_NMP_ComputeSoftmaxExp_for_1_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000)
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_2_itm_1
      , 1'b1 , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_6_0});
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_NMP_ComputeSoftmaxExp_for_1_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a
      = {NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001};
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_16_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_16_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_sva_1,
      NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_15_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_15_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_15_sva_1,
      NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_14_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_14_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_14_sva_1,
      NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_13_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_13_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_13_sva_1,
      NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_12_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_12_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_12_sva_1,
      NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_11_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_11_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_11_sva_1,
      NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_10_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_10_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_10_sva_1,
      NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_9_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_9_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_9_sva_1,
      NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_8_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_8_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_8_sva_1,
      NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_7_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_7_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_7_sva_1,
      NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_6_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_6_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_6_sva_1,
      NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_5_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_5_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_5_sva_1,
      NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_4_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_4_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_4_sva_1,
      NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_3_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_3_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_3_sva_1,
      NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_2_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_2_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_2_sva_1,
      NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_for_1_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_for_1_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_1_sva_1,
      NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_16_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_16_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_15_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_15_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_15_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_14_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_14_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_14_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_13_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_13_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_13_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_12_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_12_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_12_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_11_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_11_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_11_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_10_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_10_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_10_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_9_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_9_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_9_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_8_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_8_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_8_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_7_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_7_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_7_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_6_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_6_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_6_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_5_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_5_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_5_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_4_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_4_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_4_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_3_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_3_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_3_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_2_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_2_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_2_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [4:0] nl_NMP_ConvertOutputToAdpfloat_1_for_1_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_1_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s
      = MUX_v_5_2_2(5'b11010, out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_1_sva_1,
      NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_rg_mantissa
      = NMP_ComputeRMSNormalize_for_1_mul_cmp_1_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_rg_mantissa
      = NMP_ComputeRMSNormalize_for_1_mul_cmp_2_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_rg_mantissa
      = NMP_ComputeRMSNormalize_for_1_mul_cmp_3_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_rg_mantissa
      = NMP_ComputeRMSNormalize_for_1_mul_cmp_4_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_rg_mantissa
      = NMP_ComputeRMSNormalize_for_1_mul_cmp_5_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_rg_mantissa
      = NMP_ComputeRMSNormalize_for_1_mul_cmp_6_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_rg_mantissa
      = NMP_ComputeRMSNormalize_for_1_mul_cmp_7_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_rg_mantissa =
      NMP_ComputeRMSNormalize_for_1_mul_cmp_8_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_rg_mantissa =
      NMP_ComputeRMSNormalize_for_1_mul_cmp_9_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_rg_mantissa =
      NMP_ComputeRMSNormalize_for_1_mul_cmp_10_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_rg_mantissa =
      NMP_ComputeRMSNormalize_for_1_mul_cmp_11_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_rg_mantissa =
      NMP_ComputeRMSNormalize_for_1_mul_cmp_12_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_rg_mantissa =
      NMP_ComputeRMSNormalize_for_1_mul_cmp_13_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_rg_mantissa =
      NMP_ComputeRMSNormalize_for_1_mul_cmp_14_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_rg_mantissa =
      NMP_ComputeRMSNormalize_for_1_mul_cmp_15_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_rg_mantissa =
      NMP_ComputeRMSNormalize_for_1_mul_cmp_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_z[55:24];
  wire [31:0] nl_NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_rg_mantissa;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_rg_mantissa
      = NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_z[55:24];
  wire [36:0] nl_operator_40_0_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_operator_40_0_false_AC_TRN_AC_WRAP_lshift_rg_a = {NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_2_36_27
      , NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_2_26_0};
  wire [39:0] nl_leading_sign_40_0_rg_mantissa;
  assign nl_leading_sign_40_0_rg_mantissa = {3'b000 , NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_36_27
      , NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_26_0};
  wire[34:0] operator_40_0_false_AC_TRN_AC_WRAP_1_mux_nl;
  wire[3:0] operator_40_0_false_AC_TRN_AC_WRAP_1_operator_40_0_false_AC_TRN_AC_WRAP_1_and_nl;
  wire not_1178_nl;
  wire [38:0] nl_operator_40_0_false_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign operator_40_0_false_AC_TRN_AC_WRAP_1_mux_nl = MUX_v_35_2_2((operator_40_0_false_AC_TRN_AC_WRAP_1_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_38_0_itm[38:4]),
      sum_exp_39_4_sva_3_34_0, and_dcpl_887);
  assign not_1178_nl = ~ and_dcpl_887;
  assign operator_40_0_false_AC_TRN_AC_WRAP_1_operator_40_0_false_AC_TRN_AC_WRAP_1_and_nl
      = MUX_v_4_2_2(4'b0000, (operator_40_0_false_AC_TRN_AC_WRAP_1_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_38_0_itm[3:0]),
      not_1178_nl);
  assign nl_operator_40_0_false_AC_TRN_AC_WRAP_1_lshift_rg_a = {operator_40_0_false_AC_TRN_AC_WRAP_1_mux_nl
      , operator_40_0_false_AC_TRN_AC_WRAP_1_operator_40_0_false_AC_TRN_AC_WRAP_1_and_nl};
  wire ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_mux_nl;
  wire[34:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_mux_2_nl;
  wire[3:0] ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_and_nl;
  wire not_1179_nl;
  wire [39:0] nl_leading_sign_40_0_1_rg_mantissa;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_mux_nl
      = MUX_s_1_2_2(ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_39,
      (sum_exp_39_4_sva_2[35]), and_dcpl_893);
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_mux_2_nl
      = MUX_v_35_2_2((ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_38_0[38:4]),
      (sum_exp_39_4_sva_2[34:0]), and_dcpl_893);
  assign not_1179_nl = ~ and_dcpl_893;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_and_nl
      = MUX_v_4_2_2(4'b0000, (ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_38_0[3:0]),
      not_1179_nl);
  assign nl_leading_sign_40_0_1_rg_mantissa = {ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_mux_nl
      , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_mux_2_nl
      , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_leading_1_leading_sign_40_0_rtn_and_nl};
  wire  nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_is_write_rsc_dat_NMPRun;
  assign nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_is_write_rsc_dat_NMPRun
      = ~ NMP_RunFSM_switch_lp_conc_itm_17_0;
  wire [1:0] nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_memory_index_rsc_dat_NMPRun;
  assign nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_memory_index_rsc_dat_NMPRun
      = MUX_v_2_2_2(NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_17,
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_17, and_dcpl_581);
  wire NMP_PrepareReadReq_mux_1_nl;
  wire NMP_PrepareReadReq_mux_28_nl;
  wire[5:0] NMP_PrepareReadReq_mux_29_nl;
  wire [7:0] nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_vector_index_rsc_dat_NMPRun;
  assign NMP_PrepareReadReq_mux_1_nl = MUX_s_1_2_2(reg_NMP_PrepareReadReq_asn_1_itm_16_ftd,
      reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd, and_dcpl_581);
  assign NMP_PrepareReadReq_mux_28_nl = MUX_s_1_2_2(reg_NMP_PrepareReadReq_asn_1_itm_16_ftd_1,
      reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd_1_6, and_dcpl_581);
  assign NMP_PrepareReadReq_mux_29_nl = MUX_v_6_2_2(NMP_PrepareReadReq_asn_1_itm_16_rsp_1,
      reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd_1_5_0, and_dcpl_581);
  assign nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_vector_index_rsc_dat_NMPRun
      = {NMP_PrepareReadReq_mux_1_nl , NMP_PrepareReadReq_mux_28_nl , NMP_PrepareReadReq_mux_29_nl};
  wire[5:0] NMP_PrepareReadReq_mux_nl;
  wire[2:0] NMP_PrepareReadReq_mux_31_nl;
  wire[6:0] NMP_PrepareReadReq_mux_30_nl;
  wire [15:0] nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_timestep_index_rsc_dat_NMPRun;
  assign NMP_PrepareReadReq_mux_nl = MUX_v_6_2_2(reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_8_3,
      (reg_NMP_PrepareWriteReq_asn_2_itm_16_ftd[8:3]), and_dcpl_581);
  assign NMP_PrepareReadReq_mux_31_nl = MUX_v_3_2_2(reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_2_0,
      (reg_NMP_PrepareWriteReq_asn_2_itm_16_ftd[2:0]), and_dcpl_581);
  assign NMP_PrepareReadReq_mux_30_nl = MUX_v_7_2_2(reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_1,
      reg_NMP_PrepareWriteReq_asn_2_itm_16_ftd_1, and_dcpl_581);
  assign nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_timestep_index_rsc_dat_NMPRun
      = {NMP_PrepareReadReq_mux_nl , NMP_PrepareReadReq_mux_31_nl , NMP_PrepareReadReq_mux_30_nl};
  wire large_req_reg_write_data_data_mux_63_nl;
  wire[1:0] large_req_reg_write_data_data_mux_31_nl;
  wire large_req_reg_write_data_data_mux_30_nl;
  wire[3:0] large_req_reg_write_data_data_mux_62_nl;
  wire large_req_reg_write_data_data_mux_61_nl;
  wire[1:0] large_req_reg_write_data_data_mux_29_nl;
  wire large_req_reg_write_data_data_mux_28_nl;
  wire[3:0] large_req_reg_write_data_data_mux_60_nl;
  wire large_req_reg_write_data_data_mux_59_nl;
  wire[1:0] large_req_reg_write_data_data_mux_27_nl;
  wire large_req_reg_write_data_data_mux_26_nl;
  wire[3:0] large_req_reg_write_data_data_mux_58_nl;
  wire large_req_reg_write_data_data_mux_57_nl;
  wire[1:0] large_req_reg_write_data_data_mux_25_nl;
  wire large_req_reg_write_data_data_mux_24_nl;
  wire[3:0] large_req_reg_write_data_data_mux_56_nl;
  wire large_req_reg_write_data_data_mux_55_nl;
  wire[1:0] large_req_reg_write_data_data_mux_23_nl;
  wire large_req_reg_write_data_data_mux_22_nl;
  wire[3:0] large_req_reg_write_data_data_mux_54_nl;
  wire large_req_reg_write_data_data_mux_53_nl;
  wire[1:0] large_req_reg_write_data_data_mux_21_nl;
  wire large_req_reg_write_data_data_mux_20_nl;
  wire[3:0] large_req_reg_write_data_data_mux_52_nl;
  wire large_req_reg_write_data_data_mux_51_nl;
  wire[1:0] large_req_reg_write_data_data_mux_19_nl;
  wire large_req_reg_write_data_data_mux_18_nl;
  wire[3:0] large_req_reg_write_data_data_mux_50_nl;
  wire large_req_reg_write_data_data_mux_49_nl;
  wire[1:0] large_req_reg_write_data_data_mux_17_nl;
  wire large_req_reg_write_data_data_mux_16_nl;
  wire[3:0] large_req_reg_write_data_data_mux_48_nl;
  wire large_req_reg_write_data_data_mux_47_nl;
  wire[1:0] large_req_reg_write_data_data_mux_15_nl;
  wire large_req_reg_write_data_data_mux_14_nl;
  wire[3:0] large_req_reg_write_data_data_mux_46_nl;
  wire large_req_reg_write_data_data_mux_45_nl;
  wire[1:0] large_req_reg_write_data_data_mux_13_nl;
  wire large_req_reg_write_data_data_mux_12_nl;
  wire[3:0] large_req_reg_write_data_data_mux_44_nl;
  wire large_req_reg_write_data_data_mux_43_nl;
  wire[1:0] large_req_reg_write_data_data_mux_11_nl;
  wire large_req_reg_write_data_data_mux_10_nl;
  wire[3:0] large_req_reg_write_data_data_mux_42_nl;
  wire large_req_reg_write_data_data_mux_41_nl;
  wire[1:0] large_req_reg_write_data_data_mux_9_nl;
  wire large_req_reg_write_data_data_mux_8_nl;
  wire[3:0] large_req_reg_write_data_data_mux_40_nl;
  wire large_req_reg_write_data_data_mux_39_nl;
  wire[1:0] large_req_reg_write_data_data_mux_7_nl;
  wire large_req_reg_write_data_data_mux_6_nl;
  wire[3:0] large_req_reg_write_data_data_mux_38_nl;
  wire large_req_reg_write_data_data_mux_37_nl;
  wire[1:0] large_req_reg_write_data_data_mux_5_nl;
  wire large_req_reg_write_data_data_mux_4_nl;
  wire[3:0] large_req_reg_write_data_data_mux_36_nl;
  wire large_req_reg_write_data_data_mux_35_nl;
  wire[1:0] large_req_reg_write_data_data_mux_3_nl;
  wire large_req_reg_write_data_data_mux_2_nl;
  wire[3:0] large_req_reg_write_data_data_mux_34_nl;
  wire large_req_reg_write_data_data_mux_33_nl;
  wire[1:0] large_req_reg_write_data_data_mux_1_nl;
  wire large_req_reg_write_data_data_mux_nl;
  wire[3:0] large_req_reg_write_data_data_mux_32_nl;
  wire [127:0] nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_write_data_data_rsc_dat_NMPRun;
  assign large_req_reg_write_data_data_mux_63_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_itm_1,
      write_data_data_15_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_31_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_1_itm_1_2_1,
      write_data_data_15_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_30_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_1_itm_1_0,
      write_data_data_15_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_62_nl = MUX_v_4_2_2(large_req_reg_write_data_data_123_120_sva,
      write_data_data_15_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_61_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_3_itm_1,
      write_data_data_14_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_29_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_4_itm_1_2_1,
      write_data_data_14_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_28_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_4_itm_1_0,
      write_data_data_14_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_60_nl = MUX_v_4_2_2(large_req_reg_write_data_data_115_112_sva,
      write_data_data_14_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_59_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_6_itm_1,
      write_data_data_13_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_27_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_7_itm_1_2_1,
      write_data_data_13_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_26_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_7_itm_1_0,
      write_data_data_13_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_58_nl = MUX_v_4_2_2(large_req_reg_write_data_data_107_104_sva,
      write_data_data_13_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_57_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_9_itm_1,
      write_data_data_12_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_25_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_10_itm_1_2_1,
      write_data_data_12_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_24_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_10_itm_1_0,
      write_data_data_12_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_56_nl = MUX_v_4_2_2(large_req_reg_write_data_data_99_96_sva,
      write_data_data_12_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_55_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_12_itm_1,
      write_data_data_11_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_23_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_13_itm_1_2_1,
      write_data_data_11_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_22_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_13_itm_1_0,
      write_data_data_11_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_54_nl = MUX_v_4_2_2(large_req_reg_write_data_data_91_88_sva,
      write_data_data_11_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_53_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_15_itm_1,
      write_data_data_10_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_21_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_16_itm_1_2_1,
      write_data_data_10_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_20_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_16_itm_1_0,
      write_data_data_10_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_52_nl = MUX_v_4_2_2(large_req_reg_write_data_data_83_80_sva,
      write_data_data_10_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_51_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_18_itm_1,
      write_data_data_9_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_19_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_19_itm_1_2_1,
      write_data_data_9_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_18_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_19_itm_1_0,
      write_data_data_9_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_50_nl = MUX_v_4_2_2(large_req_reg_write_data_data_75_72_sva,
      write_data_data_9_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_49_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_21_itm_1,
      write_data_data_8_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_17_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_22_itm_1_2_1,
      write_data_data_8_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_16_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_22_itm_1_0,
      write_data_data_8_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_48_nl = MUX_v_4_2_2(large_req_reg_write_data_data_67_64_sva,
      write_data_data_8_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_47_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_24_itm_1,
      write_data_data_7_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_15_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_25_itm_1_2_1,
      write_data_data_7_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_14_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_25_itm_1_0,
      write_data_data_7_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_46_nl = MUX_v_4_2_2(large_req_reg_write_data_data_59_56_sva,
      write_data_data_7_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_45_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_27_itm_1,
      write_data_data_6_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_13_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_28_itm_1_2_1,
      write_data_data_6_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_12_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_28_itm_1_0,
      write_data_data_6_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_44_nl = MUX_v_4_2_2(large_req_reg_write_data_data_51_48_sva,
      write_data_data_6_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_43_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_30_itm_1,
      write_data_data_5_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_11_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_31_itm_1_2_1,
      write_data_data_5_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_10_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_31_itm_1_0,
      write_data_data_5_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_42_nl = MUX_v_4_2_2(large_req_reg_write_data_data_43_40_sva,
      write_data_data_5_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_41_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_33_itm_1,
      write_data_data_4_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_9_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_34_itm_1_2_1,
      write_data_data_4_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_8_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_34_itm_1_0,
      write_data_data_4_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_40_nl = MUX_v_4_2_2(large_req_reg_write_data_data_35_32_sva,
      write_data_data_4_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_39_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_36_itm_1,
      write_data_data_3_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_7_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_37_itm_1_2_1,
      write_data_data_3_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_6_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_37_itm_1_0,
      write_data_data_3_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_38_nl = MUX_v_4_2_2(large_req_reg_write_data_data_27_24_sva,
      write_data_data_3_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_37_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_39_itm_1,
      write_data_data_2_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_5_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_40_itm_1_2_1,
      write_data_data_2_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_4_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_40_itm_1_0,
      write_data_data_2_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_36_nl = MUX_v_4_2_2(large_req_reg_write_data_data_19_16_sva,
      write_data_data_2_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_35_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_42_itm_1,
      write_data_data_1_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_3_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_43_itm_1_2_1,
      write_data_data_1_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_2_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_43_itm_1_0,
      write_data_data_1_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_34_nl = MUX_v_4_2_2(large_req_reg_write_data_data_11_8_sva,
      write_data_data_1_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_33_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_45_itm_1,
      write_data_data_0_7_sva_dfm_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_1_nl = MUX_v_2_2_2(large_req_reg_write_data_data_asn_46_itm_1_2_1,
      write_data_data_0_6_4_sva_dfm_1_2_1, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_nl = MUX_s_1_2_2(large_req_reg_write_data_data_asn_46_itm_1_0,
      write_data_data_0_6_4_sva_dfm_1_0, and_dcpl_581);
  assign large_req_reg_write_data_data_mux_32_nl = MUX_v_4_2_2(large_req_reg_write_data_data_3_0_sva,
      write_data_data_0_3_0_sva_dfm_1_mx1, and_dcpl_581);
  assign nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_write_data_data_rsc_dat_NMPRun
      = {large_req_reg_write_data_data_mux_63_nl , large_req_reg_write_data_data_mux_31_nl
      , large_req_reg_write_data_data_mux_30_nl , large_req_reg_write_data_data_mux_62_nl
      , large_req_reg_write_data_data_mux_61_nl , large_req_reg_write_data_data_mux_29_nl
      , large_req_reg_write_data_data_mux_28_nl , large_req_reg_write_data_data_mux_60_nl
      , large_req_reg_write_data_data_mux_59_nl , large_req_reg_write_data_data_mux_27_nl
      , large_req_reg_write_data_data_mux_26_nl , large_req_reg_write_data_data_mux_58_nl
      , large_req_reg_write_data_data_mux_57_nl , large_req_reg_write_data_data_mux_25_nl
      , large_req_reg_write_data_data_mux_24_nl , large_req_reg_write_data_data_mux_56_nl
      , large_req_reg_write_data_data_mux_55_nl , large_req_reg_write_data_data_mux_23_nl
      , large_req_reg_write_data_data_mux_22_nl , large_req_reg_write_data_data_mux_54_nl
      , large_req_reg_write_data_data_mux_53_nl , large_req_reg_write_data_data_mux_21_nl
      , large_req_reg_write_data_data_mux_20_nl , large_req_reg_write_data_data_mux_52_nl
      , large_req_reg_write_data_data_mux_51_nl , large_req_reg_write_data_data_mux_19_nl
      , large_req_reg_write_data_data_mux_18_nl , large_req_reg_write_data_data_mux_50_nl
      , large_req_reg_write_data_data_mux_49_nl , large_req_reg_write_data_data_mux_17_nl
      , large_req_reg_write_data_data_mux_16_nl , large_req_reg_write_data_data_mux_48_nl
      , large_req_reg_write_data_data_mux_47_nl , large_req_reg_write_data_data_mux_15_nl
      , large_req_reg_write_data_data_mux_14_nl , large_req_reg_write_data_data_mux_46_nl
      , large_req_reg_write_data_data_mux_45_nl , large_req_reg_write_data_data_mux_13_nl
      , large_req_reg_write_data_data_mux_12_nl , large_req_reg_write_data_data_mux_44_nl
      , large_req_reg_write_data_data_mux_43_nl , large_req_reg_write_data_data_mux_11_nl
      , large_req_reg_write_data_data_mux_10_nl , large_req_reg_write_data_data_mux_42_nl
      , large_req_reg_write_data_data_mux_41_nl , large_req_reg_write_data_data_mux_9_nl
      , large_req_reg_write_data_data_mux_8_nl , large_req_reg_write_data_data_mux_40_nl
      , large_req_reg_write_data_data_mux_39_nl , large_req_reg_write_data_data_mux_7_nl
      , large_req_reg_write_data_data_mux_6_nl , large_req_reg_write_data_data_mux_38_nl
      , large_req_reg_write_data_data_mux_37_nl , large_req_reg_write_data_data_mux_5_nl
      , large_req_reg_write_data_data_mux_4_nl , large_req_reg_write_data_data_mux_36_nl
      , large_req_reg_write_data_data_mux_35_nl , large_req_reg_write_data_data_mux_3_nl
      , large_req_reg_write_data_data_mux_2_nl , large_req_reg_write_data_data_mux_34_nl
      , large_req_reg_write_data_data_mux_33_nl , large_req_reg_write_data_data_mux_1_nl
      , large_req_reg_write_data_data_mux_nl , large_req_reg_write_data_data_mux_32_nl};
  wire [127:0] nl_NMP_NMPRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff;
  assign nl_NMP_NMPRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff
      = {29'b00000000000000000000000000000 , rva_out_reg_data_98_96_sva_dfm_3_17_2
      , rva_out_reg_data_98_96_sva_dfm_3_17_1_0 , 16'b0000000000000000 , rva_out_reg_data_79_64_sva_dfm_3_17
      , 8'b00000000 , rva_out_reg_data_55_48_sva_dfm_3_17 , 13'b0000000000000 , rva_out_reg_data_34_32_sva_dfm_3_17
      , 21'b000000000000000000000 , rva_out_reg_data_10_8_sva_dfm_3_17 , 7'b0000000
      , rva_out_reg_data_0_sva_dfm_3_17};
  GBModule_mgc_shift_br_v5 #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_s(32'sd7),
  .width_z(32'sd40)) operator_40_16_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_operator_40_16_true_AC_TRN_AC_WRAP_rshift_rg_a[25:0]),
      .s(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_3),
      .z(operator_40_16_true_AC_TRN_AC_WRAP_rshift_itm)
    );
  GBModule_mgc_shift_br_v5 #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd40)) operator_40_16_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_operator_40_16_true_AC_TRN_AC_WRAP_1_rshift_rg_a[24:0]),
      .s(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_3),
      .z(operator_40_16_true_AC_TRN_AC_WRAP_1_rshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd27)) NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_rg
      (
      .a(nl_NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_rg_a[21:0]),
      .s(nl_NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_rg_s[4:0]),
      .z(NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd40)) operator_40_16_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_40_16_false_AC_TRN_AC_WRAP_lshift_rg_a[24:0]),
      .s(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_6_1_itm_1),
      .z(operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_16_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_16_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_16_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_16_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_15_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_15_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_15_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_15_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_14_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_14_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_14_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_14_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_13_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_13_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_13_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_13_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_12_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_12_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_12_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_12_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_11_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_11_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_11_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_11_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_10_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_10_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_8_0),
      .z(NMP_ComputeSoftmaxExp_for_10_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_9_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_9_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_9_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_9_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_8_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_8_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_8_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_8_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_7_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_7_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_7_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_7_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_6_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_6_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_6_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_6_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_5_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_5_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_5_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_5_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_4_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_4_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_4_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_4_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_3_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_3_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_3_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_3_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_2_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_2_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_2_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_2_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd32)) NMP_ComputeSoftmaxExp_for_1_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(nl_NMP_ComputeSoftmaxExp_for_1_operator_32_12_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1),
      .z(NMP_ComputeSoftmaxExp_for_1_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_16_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_16_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_16_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_16_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_15_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_15_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_15_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_15_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_14_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_14_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_14_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_14_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_13_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_13_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_13_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_13_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_12_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_12_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_12_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_12_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_11_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_11_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_11_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_11_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_10_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_10_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_10_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_10_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_9_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_9_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_9_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_9_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_8_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_8_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_8_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_8_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_7_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_7_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_7_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_7_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_6_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_6_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_6_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_6_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_5_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_5_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_5_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_5_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_4_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_4_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_4_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_4_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_3_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_3_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_3_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_3_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_2_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_2_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_2_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_2_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_for_1_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg
      (
      .a(NMP_ComputeRMSNormalize_for_1_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_for_1_operator_32_12_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_for_1_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_16_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_16_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_16_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_16_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_15_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_15_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_15_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_15_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_14_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_14_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_14_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_14_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_13_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_13_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_13_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_13_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_12_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_12_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_12_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_12_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_11_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_11_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_11_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_11_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_10_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_10_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_10_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_10_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_9_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_9_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_9_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_9_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_8_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_8_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_8_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_8_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_7_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_7_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_7_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_7_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_6_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_6_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_6_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_6_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_5_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_5_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_5_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_5_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_4_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_4_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_4_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_4_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_3_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_3_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_3_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_3_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_2_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_2_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_2_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_2_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd32)) NMP_ConvertOutputToAdpfloat_1_for_1_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg
      (
      .a(NMP_ComputeSoftmaxNormalize_for_1_slc_55_24_ncse_sva_1),
      .s(nl_NMP_ConvertOutputToAdpfloat_1_for_1_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(NMP_ConvertOutputToAdpfloat_1_for_1_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_leading_sign_32_1_1_0  NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_rg
      (
      .mantissa(nl_NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_rg_mantissa[31:0]),
      .all_same(NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_out_2),
      .rtn(NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_out_3)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd37),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd39)) operator_40_0_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_40_0_false_AC_TRN_AC_WRAP_lshift_rg_a[36:0]),
      .s(NMP_PrepareReadReq_asn_1_itm_4_5_0),
      .z(operator_40_0_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  GBModule_leading_sign_40_0  leading_sign_40_0_rg (
      .mantissa(nl_leading_sign_40_0_rg_mantissa[39:0]),
      .rtn(leading_sign_40_0_out_1)
    );
  GBModule_mgc_shift_l_v5 #(.width_a(32'sd39),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd39)) operator_40_0_false_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_operator_40_0_false_AC_TRN_AC_WRAP_1_lshift_rg_a[38:0]),
      .s(NMP_PrepareReadReq_asn_1_itm_10_5_0),
      .z(z_out_2)
    );
  GBModule_leading_sign_40_0  leading_sign_40_0_1_rg (
      .mantissa(nl_leading_sign_40_0_1_rg_mantissa[39:0]),
      .rtn(rtn_out)
    );
  GBModule_NMP_NMPRun_rva_in_PopNB_mioi NMP_NMPRun_rva_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .NMPRun_wen(NMPRun_wen),
      .NMPRun_wten(NMPRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(fsm_output)
    );
  GBModule_NMP_NMPRun_large_req_Push_mioi NMP_NMPRun_large_req_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .large_req_vld(large_req_vld),
      .large_req_rdy(large_req_rdy),
      .large_req_dat(large_req_dat),
      .NMPRun_wen(NMPRun_wen),
      .large_req_Push_mioi_oswt(reg_large_req_Push_mioi_iswt0_cse),
      .large_req_Push_mioi_wen_comp(large_req_Push_mioi_wen_comp),
      .large_req_Push_mioi_m_is_write_rsc_dat_NMPRun(nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_is_write_rsc_dat_NMPRun),
      .large_req_Push_mioi_m_memory_index_rsc_dat_NMPRun(nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_memory_index_rsc_dat_NMPRun[1:0]),
      .large_req_Push_mioi_m_vector_index_rsc_dat_NMPRun(nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_vector_index_rsc_dat_NMPRun[7:0]),
      .large_req_Push_mioi_m_timestep_index_rsc_dat_NMPRun(nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_timestep_index_rsc_dat_NMPRun[15:0]),
      .large_req_Push_mioi_m_write_data_data_rsc_dat_NMPRun(nl_NMP_NMPRun_large_req_Push_mioi_inst_large_req_Push_mioi_m_write_data_data_rsc_dat_NMPRun[127:0]),
      .large_req_Push_mioi_oswt_pff(nor_206_rmff)
    );
  GBModule_NMP_NMPRun_start_PopNB_mioi NMP_NMPRun_start_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .NMPRun_wen(NMPRun_wen),
      .NMPRun_wten(NMPRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_oswt_pff(and_591_rmff)
    );
  GBModule_NMP_NMPRun_large_rsp_PopNB_mioi NMP_NMPRun_large_rsp_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .large_rsp_vld(large_rsp_vld),
      .large_rsp_rdy(large_rsp_rdy),
      .large_rsp_dat(large_rsp_dat),
      .NMPRun_wen(NMPRun_wen),
      .NMPRun_wten(NMPRun_wten),
      .large_rsp_PopNB_mioi_oswt(reg_large_rsp_PopNB_mioi_iswt0_cse),
      .large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt),
      .large_rsp_PopNB_mioi_return_rsc_z_mxwt(large_rsp_PopNB_mioi_return_rsc_z_mxwt),
      .large_rsp_PopNB_mioi_oswt_pff(and_590_rmff)
    );
  GBModule_NMP_NMPRun_rva_out_Push_mioi NMP_NMPRun_rva_out_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .NMPRun_wen(NMPRun_wen),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff(nl_NMP_NMPRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_NMPRun_pff[127:0]),
      .rva_out_Push_mioi_oswt_pff(and_588_rmff)
    );
  GBModule_NMP_NMPRun_done_Push_mioi NMP_NMPRun_done_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .done_vld(done_vld),
      .done_rdy(done_rdy),
      .done_dat(done_dat),
      .NMPRun_wen(NMPRun_wen),
      .done_Push_mioi_oswt(reg_done_Push_mioi_iswt0_cse),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp),
      .done_Push_mioi_oswt_pff(and_587_rmff)
    );
  GBModule_NMP_NMPRun_wait_dp NMP_NMPRun_wait_dp_inst (
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .NMPRun_wen(NMPRun_wen),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo(reg_NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo_ir_15_cse),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo_ir_unreg(and_585_rmff),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo(reg_NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo_ir_15_cse),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo_ir_unreg(and_584_rmff),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo(reg_NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo_ir_15_cse),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo_ir_unreg(and_583_rmff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo(reg_NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo_ir_15_cse),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo_ir_unreg(and_582_rmff)
    );
  GBModule_NMP_NMPRun_staller NMP_NMPRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .NMPRun_wen(NMPRun_wen),
      .NMPRun_wten(NMPRun_wten),
      .large_req_Push_mioi_wen_comp(large_req_Push_mioi_wen_comp),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp)
    );
  GBModule_NMP_NMPRun_NMPRun_fsm NMP_NMPRun_NMPRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .NMPRun_wen(NMPRun_wen),
      .fsm_output(fsm_output)
    );
  assign nor_201_nl = ~(state_0_sva | (~ or_tmp_35));
  assign or_504_nl = (~ while_stage_0_3) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ state_1_sva) | state_3_sva | state_2_sva;
  assign mux_16_nl = MUX_s_1_2_2(nor_201_nl, or_tmp_35, or_504_nl);
  assign and_582_rmff = (~ mux_16_nl) & fsm_output;
  assign nor_202_nl = ~(while_stage_0_14 | (~ mux_tmp_17));
  assign or_508_nl = (~ NMP_RunFSM_switch_lp_conc_itm_12_0) | (~ NMP_RunFSM_switch_lp_conc_itm_12_2)
      | NMP_RunFSM_switch_lp_conc_itm_12_3 | NMP_RunFSM_switch_lp_conc_itm_12_1 |
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_12;
  assign mux_18_nl = MUX_s_1_2_2(nor_202_nl, mux_tmp_17, or_508_nl);
  assign and_583_rmff = (~ mux_18_nl) & fsm_output;
  assign nor_203_nl = ~(while_stage_0_8 | (~ or_tmp_45));
  assign or_514_nl = NMP_RunFSM_switch_lp_conc_itm_6_3 | (~ NMP_RunFSM_switch_lp_conc_itm_6_2)
      | (~ NMP_RunFSM_switch_lp_conc_itm_6_0) | (~ NMP_RunFSM_switch_lp_conc_itm_6_1)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  assign mux_19_nl = MUX_s_1_2_2(nor_203_nl, or_tmp_45, or_514_nl);
  assign and_584_rmff = (~ mux_19_nl) & fsm_output;
  assign nor_204_nl = ~(while_stage_0_14 | (~ mux_tmp_20));
  assign or_518_nl = (~ NMP_RunFSM_switch_lp_conc_itm_12_0) | NMP_RunFSM_switch_lp_conc_itm_12_2
      | (~ NMP_RunFSM_switch_lp_conc_itm_12_3) | NMP_RunFSM_switch_lp_conc_itm_12_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_12;
  assign mux_21_nl = MUX_s_1_2_2(nor_204_nl, mux_tmp_20, or_518_nl);
  assign and_585_rmff = (~ mux_21_nl) & fsm_output;
  assign and_587_rmff = while_stage_0_19 & (~ while_while_nor_itm_17) & while_while_and_itm_17;
  assign and_588_rmff = while_stage_0_19 & while_while_nor_itm_17;
  assign or_533_cse = (~ NMP_RunFSM_switch_lp_or_73_tmp) | NMP_UpdateFSM_switch_lp_equal_tmp_1
      | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign or_534_cse = state_0_sva | state_3_sva;
  assign or_536_nl = (~ is_start_sva) | NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign or_535_nl = (~ start_PopNB_mioi_data_rsc_z_mxwt) | (~ nmp_config_is_valid_sva)
      | NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign mux_38_nl = MUX_s_1_2_2(or_536_nl, or_535_nl, start_PopNB_mioi_return_rsc_z_mxwt);
  assign mux_41_nl = MUX_s_1_2_2(mux_38_nl, or_803_cse, or_tmp_56);
  assign mux_45_nl = MUX_s_1_2_2(mux_tmp_25, mux_41_nl, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_46_nl = MUX_s_1_2_2(mux_45_nl, mux_tmp_26, or_534_cse);
  assign mux_24_nl = MUX_s_1_2_2(or_tmp_60, or_803_cse, next_state_3_lpi_1_dfm_3);
  assign mux_33_nl = MUX_s_1_2_2(or_tmp_60, or_803_cse, large_rsp_PopNB_mioi_return_rsc_z_mxwt);
  assign mux_34_nl = MUX_s_1_2_2(mux_24_nl, mux_33_nl, NMP_RunFSM_switch_lp_equal_tmp_11_1);
  assign nor_5_nl = ~(NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2 | (~ large_rsp_PopNB_mioi_return_rsc_z_mxwt));
  assign mux_30_nl = MUX_s_1_2_2(or_tmp_57, or_803_cse, nor_5_nl);
  assign mux_32_nl = MUX_s_1_2_2(or_tmp_57, mux_30_nl, NMP_RunFSM_switch_lp_equal_tmp_11_1);
  assign mux_35_nl = MUX_s_1_2_2(mux_34_nl, mux_32_nl, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_36_nl = MUX_s_1_2_2(mux_35_nl, mux_tmp_26, state_3_sva);
  assign mux_28_nl = MUX_s_1_2_2(mux_tmp_25, or_533_cse, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign or_532_nl = (~ state_3_sva) | nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1
      | operator_16_false_acc_2_itm_17;
  assign mux_29_nl = MUX_s_1_2_2(mux_28_nl, mux_tmp_26, or_532_nl);
  assign mux_37_nl = MUX_s_1_2_2(mux_36_nl, mux_29_nl, state_0_sva);
  assign mux_47_nl = MUX_s_1_2_2(mux_46_nl, mux_37_nl, state_1_sva);
  assign mux_48_nl = MUX_s_1_2_2(mux_47_nl, mux_tmp_26, state_2_sva);
  assign or_538_nl = NMP_UpdateFSM_switch_lp_equal_tmp_1_1 | NMP_UpdateFSM_switch_lp_equal_tmp_4_1
      | NMP_UpdateFSM_switch_lp_or_tmp_1 | NMP_UpdateFSM_switch_lp_equal_tmp_2_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_3_1 | NMP_UpdateFSM_switch_lp_equal_tmp_5_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_6_1 | (~ mux_48_nl);
  assign or_524_nl = state_2_sva | state_0_sva | state_3_sva;
  assign mux_49_cse = MUX_s_1_2_2(or_538_nl, or_524_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nor_205_nl = ~(state_2_sva | (~ state_1_sva) | state_0_sva | state_3_sva);
  assign and_893_nl = state_1_sva_dfm_1 & (~ mux_49_cse);
  assign mux_50_nl = MUX_s_1_2_2(nor_205_nl, and_893_nl, while_stage_0_3);
  assign and_590_rmff = mux_50_nl & and_dcpl_172;
  assign or_555_nl = state_1_sva_dfm_1 | mux_49_cse;
  assign mux_79_nl = MUX_s_1_2_2(or_tmp_85, or_555_nl, while_stage_0_3);
  assign and_591_rmff = (~ mux_79_nl) & and_dcpl_172;
  assign or_557_nl = (~ NMP_RunFSM_switch_lp_conc_itm_17_1) | NMP_RunFSM_switch_lp_conc_itm_17_0;
  assign mux_80_nl = MUX_s_1_2_2(or_tmp_87, or_557_nl, NMP_RunFSM_switch_lp_conc_itm_17_3);
  assign nor_206_rmff = ~(mux_80_nl | (~ while_stage_0_19) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17
      | NMP_RunFSM_switch_lp_conc_itm_17_2);
  assign or_928_cse = NMP_RunFSM_switch_lp_equal_tmp_13_1 | NMP_RunFSM_switch_lp_equal_tmp_3_12;
  assign NMP_RunFSM_switch_lp_and_7_nl = ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_4
      & NMP_RunFSM_switch_lp_equal_tmp_3_12;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux_nl =
      MUX_v_40_2_2(40'b0111111111111111111111111111111111111111, operator_40_16_true_AC_TRN_AC_WRAP_rshift_itm,
      NMP_RunFSM_switch_lp_and_7_nl);
  assign NMP_RunFSM_switch_lp_not_63_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_13_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_33_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux_nl, NMP_RunFSM_switch_lp_not_63_nl);
  assign rms_reciprocal_and_nl = or_928_cse & and_dcpl_97 & fsm_output;
  assign rms_reciprocal_mux_rmff = MUX_v_40_2_2(reg_NMP_ComputeRMSNormalize_for_1_mul_cmp_15_b_cse,
      NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_33_nl, rms_reciprocal_and_nl);
  assign or_929_cse = NMP_RunFSM_switch_lp_equal_tmp_13_1 | NMP_RunFSM_switch_lp_equal_tmp_7_12;
  assign NMP_RunFSM_switch_lp_and_5_nl = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_5
      & NMP_RunFSM_switch_lp_equal_tmp_7_12;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux_1_nl
      = MUX_v_40_2_2(40'b0111111111111111111111111111111111111111, operator_40_16_true_AC_TRN_AC_WRAP_1_rshift_itm,
      NMP_RunFSM_switch_lp_and_5_nl);
  assign NMP_RunFSM_switch_lp_not_49_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_13_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_32_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux_1_nl, NMP_RunFSM_switch_lp_not_49_nl);
  assign sum_exp_reciprocal_and_nl = or_929_cse & and_dcpl_97 & fsm_output;
  assign sum_exp_reciprocal_mux_rmff = MUX_v_40_2_2(reg_NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_b_cse,
      NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_32_nl, sum_exp_reciprocal_and_nl);
  assign and_936_cse = (NMP_RunFSM_switch_lp_equal_tmp_4_17 | NMP_RunFSM_switch_lp_equal_tmp_8_17)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_18)
      & NMPRun_wen & while_stage_0_20;
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse = NMPRun_wen & and_dcpl
      & NMP_RunFSM_switch_lp_equal_tmp_4_16;
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_16_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_15_itm_1_enexo
      | reg_out_float_round_32_if_m_1_1_sva_1_3_0_enexo | reg_out_float_round_32_if_m_1_1_sva_1_6_enexo
      | reg_NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse = NMPRun_wen & and_dcpl
      & NMP_RunFSM_switch_lp_equal_tmp_8_16;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_16_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_15_itm_1_enexo
      | reg_NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_1_sva_1_3_0_enexo | reg_out_float_round_32_1_if_m_1_1_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_17_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1_enexo
      | reg_out_float_round_32_if_m_1_17_sva_1_3_0_enexo | reg_out_float_round_32_if_m_1_17_sva_1_6_enexo
      | reg_NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_17_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_14_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_17_sva_1_6_enexo | reg_NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_17_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_18_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_13_itm_1_enexo
      | reg_out_float_round_32_if_m_1_16_sva_1_3_0_enexo | reg_NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
      | reg_out_float_round_32_if_m_1_16_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_18_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_16_sva_1_3_0_enexo | reg_NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_16_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_19_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_out_float_round_32_if_m_1_15_sva_1_3_0_enexo | reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_3
      | reg_out_float_round_32_if_m_1_15_sva_1_6_enexo | reg_NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_19_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_12_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_15_sva_1_6_enexo | reg_out_float_round_32_1_if_m_1_15_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_20_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1_enexo
      | reg_out_float_round_32_if_m_1_14_sva_1_6_enexo | reg_out_float_round_32_if_m_1_14_sva_1_3_0_enexo
      | reg_NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_20_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_11_itm_1_enexo
      | reg_NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_14_sva_1_3_0_enexo | reg_out_float_round_32_1_if_m_1_14_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_21_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1_enexo
      | reg_NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
      | reg_out_float_round_32_if_m_1_13_sva_1_6_enexo | reg_out_float_round_32_if_m_1_13_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_21_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_10_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_13_sva_1_6_enexo | reg_NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_13_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_22_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
      | reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1_enexo
      | reg_out_float_round_32_if_m_1_12_sva_1_6_enexo | reg_out_float_round_32_if_m_1_12_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_22_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1_enexo
      | reg_NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_12_sva_1_6_enexo | reg_out_float_round_32_1_if_m_1_12_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_23_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_7 | reg_NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
      | reg_out_float_round_32_if_m_1_11_sva_1_3_0_enexo | reg_out_float_round_32_if_m_1_11_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_23_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_8_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_11_sva_1_6_enexo | reg_NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_11_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_24_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1_enexo
      | reg_out_float_round_32_if_m_1_10_sva_1_6_enexo | reg_out_float_round_32_if_m_1_10_sva_1_3_0_enexo
      | reg_NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_24_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_10_sva_1_3_0_enexo | reg_NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_10_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_25_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_out_float_round_32_if_m_1_9_sva_1_3_0_enexo | reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_6_itm_1_enexo
      | reg_out_float_round_32_if_m_1_9_sva_1_6_enexo | reg_NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_25_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_out_float_round_32_1_if_m_1_9_sva_1_6_enexo | reg_NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_9_sva_1_3_0_enexo | reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_6_itm_1_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_26_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1_enexo
      | reg_out_float_round_32_if_m_1_8_sva_1_6_enexo | reg_NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
      | reg_out_float_round_32_if_m_1_8_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_26_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_8_sva_1_3_0_enexo | reg_out_float_round_32_1_if_m_1_8_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_27_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1_enexo
      | reg_out_float_round_32_if_m_1_7_sva_1_3_0_enexo | reg_out_float_round_32_if_m_1_7_sva_1_6_enexo
      | reg_NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_27_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_4_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_7_sva_1_6_enexo | reg_out_float_round_32_1_if_m_1_7_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_28_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_out_float_round_32_if_m_1_6_sva_1_6_enexo | reg_out_float_round_32_if_m_1_6_sva_1_3_0_enexo
      | reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_3_itm_1_enexo
      | reg_NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_28_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_out_float_round_32_1_if_m_1_6_sva_1_3_0_enexo | reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1_enexo
      | reg_NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_6_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_29_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
      | reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_2_itm_1_enexo
      | reg_out_float_round_32_if_m_1_5_sva_1_6_enexo | reg_out_float_round_32_if_m_1_5_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_29_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_5_sva_1_3_0_enexo | reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_5_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_30_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_14 | reg_NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
      | reg_out_float_round_32_if_m_1_4_sva_1_3_0_enexo | reg_out_float_round_32_if_m_1_4_sva_1_6_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_30_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_4_sva_1_6_enexo | reg_NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_out_float_round_32_1_if_m_1_4_sva_1_3_0_enexo);
  assign NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_31_enex5 = NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_cse
      & (reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_itm_1_enexo
      | reg_out_float_round_32_if_m_1_3_sva_1_6_enexo | reg_out_float_round_32_if_m_1_3_sva_1_3_0_enexo
      | reg_NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_31_enex5 = NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_cse
      & (reg_out_float_round_32_1_if_m_1_3_sva_1_3_0_enexo | reg_NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
      | reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1_enexo
      | reg_out_float_round_32_1_if_m_1_3_sva_1_6_enexo);
  assign NMP_RunFSM_switch_lp_and_cse = NMPRun_wen & while_stage_0_19;
  assign large_req_reg_write_data_data_and_64_cse = NMPRun_wen & and_dcpl_6 & and_dcpl_3
      & (~ NMP_RunFSM_switch_lp_conc_itm_16_3);
  assign large_req_reg_write_data_data_and_cse = NMPRun_wen & (~(or_dcpl_471 | (~
      NMP_RunFSM_switch_lp_equal_tmp_9_16)));
  assign NMP_PrepareReadReq_and_55_enex5 = large_req_reg_write_data_data_and_64_cse
      & reg_NMP_PrepareReadReq_asn_2_itm_15_1_enexo;
  assign in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse = NMPRun_wen & and_dcpl_6
      & NMP_RunFSM_switch_lp_conc_itm_16_0 & NMP_RunFSM_switch_lp_conc_itm_16_2 &
      (~ NMP_RunFSM_switch_lp_conc_itm_16_3);
  assign in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse = NMPRun_wen & and_dcpl_6
      & and_dcpl_3 & NMP_RunFSM_switch_lp_conc_itm_16_3;
  assign write_data_data_and_16_cse = NMPRun_wen & (~ or_dcpl_471);
  assign NMP_PrepareWriteReq_and_12_cse = NMPRun_wen & and_dcpl_5 & NMP_RunFSM_switch_lp_conc_itm_16_1
      & (~(NMP_RunFSM_switch_lp_conc_itm_16_0 | NMP_RunFSM_switch_lp_conc_itm_16_2))
      & NMP_RunFSM_switch_lp_conc_itm_16_3;
  assign NMP_PrepareWriteReq_and_61_enex5 = NMP_PrepareWriteReq_and_12_cse & reg_NMP_PrepareWriteReq_asn_2_itm_15_enexo;
  assign NMP_PrepareWriteReq_and_62_enex5 = NMP_PrepareWriteReq_and_12_cse & reg_NMP_PrepareWriteReq_asn_2_itm_15_1_enexo;
  assign NMP_RunFSM_switch_lp_and_39_cse = NMPRun_wen & and_dcpl_5;
  assign rva_out_reg_data_and_6_cse = NMPRun_wen & while_while_nor_itm_16 & while_stage_0_18;
  assign rva_out_reg_data_and_102_enex5 = rva_out_reg_data_and_6_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_16_enexo;
  assign rva_out_reg_data_and_103_enex5 = rva_out_reg_data_and_6_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_16_enexo;
  assign while_and_144_cse = NMPRun_wen & while_stage_0_18;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_cse = NMPRun_wen &
      and_dcpl_91 & and_dcpl_88 & NMP_RunFSM_switch_lp_conc_itm_15_2;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_cse = NMPRun_wen
      & and_dcpl_91 & (~ NMP_RunFSM_switch_lp_conc_itm_15_1) & NMP_RunFSM_switch_lp_conc_itm_15_3
      & (~ NMP_RunFSM_switch_lp_conc_itm_15_2);
  assign NMP_RunFSM_switch_lp_and_43_cse = NMPRun_wen & and_dcpl_90;
  assign while_if_and_2_cse = NMPRun_wen & while_stage_0_17;
  assign NMP_RunFSM_switch_lp_and_47_cse = NMPRun_wen & and_dcpl_96;
  assign while_if_and_3_cse = NMPRun_wen & while_stage_0_16;
  assign NMP_RunFSM_switch_lp_and_51_cse = NMPRun_wen & and_dcpl_97;
  assign while_if_and_4_cse = NMPRun_wen & while_stage_0_15;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5
      = NMPRun_wen & (reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_3_enexo
      | reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_enexo);
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_3_enex5 = NMPRun_wen
      & reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_2_enexo;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_1_enex5
      = NMPRun_wen & ((sum_exp_39_4_sva_st_4!=36'b000000000000000000000000000000000000))
      & and_dcpl_108 & NMP_RunFSM_switch_lp_equal_tmp_7_11 & (~ NMP_RunFSM_switch_lp_conc_itm_12_1)
      & and_dcpl_105 & (~ NMP_RunFSM_switch_lp_conc_itm_12_0) & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_4
      & reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_2_enexo;
  assign NMP_RunFSM_switch_lp_and_55_cse = NMPRun_wen & while_stage_0_14;
  assign NMP_RunFSM_switch_lp_and_56_cse = NMPRun_wen & and_dcpl_108;
  assign NMP_RunFSM_switch_lp_and_60_cse = NMPRun_wen & and_dcpl_100;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_enex5
      = NMPRun_wen & and_dcpl_125 & and_dcpl_122 & (~ NMP_RunFSM_switch_lp_conc_itm_11_0)
      & reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_2_enexo;
  assign NMP_ComputeRMSNormalize_for_and_cse = NMPRun_wen & and_dcpl_125 & and_dcpl_122
      & NMP_RunFSM_switch_lp_conc_itm_11_0;
  assign NMP_ComputeRMSNormalize_for_and_145_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_60_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_146_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_58_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_147_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_56_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_148_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_54_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_149_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_52_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_150_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_50_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_151_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_48_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_152_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_46_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_153_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_44_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_154_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_42_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_155_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_40_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_156_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_38_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_157_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_36_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_158_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_34_itm_10_enexo;
  assign NMP_ComputeRMSNormalize_for_and_159_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_32_itm_10_enexo;
  assign NMP_ComputeRMSNormalize_for_and_160_enex5 = NMP_ComputeRMSNormalize_for_and_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_itm_10_enexo;
  assign sum_exp_and_enex5 = NMPRun_wen & and_dcpl_125 & and_dcpl_130 & reg_sum_exp_39_4_sva_st_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_cse = NMPRun_wen & and_dcpl_125 & and_dcpl_129
      & NMP_RunFSM_switch_lp_conc_itm_11_0;
  assign NMP_ComputeSoftmaxNormalize_for_and_80_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_81_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_82_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_83_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_84_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_85_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_86_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_87_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_88_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_89_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_90_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_91_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_92_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_93_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_94_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_95_enex5 = NMP_ComputeSoftmaxNormalize_for_and_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_3_enexo;
  assign NMP_RunFSM_switch_lp_and_64_cse = NMPRun_wen & and_dcpl_124;
  assign while_if_and_6_cse = NMPRun_wen & while_stage_0_13;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_1_enex5
      = NMPRun_wen & and_dcpl_137 & and_dcpl_134 & (~ NMP_RunFSM_switch_lp_conc_itm_10_0)
      & reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_1_enexo;
  assign sum_exp_and_1_enex5 = NMPRun_wen & and_dcpl_142 & reg_sum_exp_39_4_sva_st_2_enexo;
  assign NMP_RunFSM_switch_lp_and_68_cse = NMPRun_wen & and_dcpl_136;
  assign while_if_and_7_cse = NMPRun_wen & while_stage_0_12;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_2_cse
      = NMPRun_wen & and_dcpl_146 & and_dcpl_143 & (~ NMP_RunFSM_switch_lp_conc_itm_9_0);
  assign sum_exp_and_2_enex5 = NMPRun_wen & and_dcpl_150 & and_dcpl_148 & (~ NMP_RunFSM_switch_lp_conc_itm_9_0)
      & reg_sum_exp_39_4_sva_st_1_enexo;
  assign NMP_RunFSM_switch_lp_and_72_cse = NMPRun_wen & and_dcpl_145;
  assign while_if_and_8_cse = NMPRun_wen & while_stage_0_11;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_2_cse
      = NMPRun_wen & and_dcpl_155 & and_dcpl_152 & (~ NMP_RunFSM_switch_lp_conc_itm_8_0);
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_12_enex5 = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_2_cse
      & reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo;
  assign NMP_RunFSM_switch_lp_and_76_cse = NMPRun_wen & and_dcpl_154;
  assign while_if_and_9_cse = NMPRun_wen & while_stage_0_10;
  assign NMP_RunFSM_switch_lp_and_80_cse = NMPRun_wen & and_dcpl_159;
  assign while_if_and_10_cse = NMPRun_wen & while_stage_0_9;
  assign NMP_RunFSM_switch_lp_and_84_cse = NMPRun_wen & and_dcpl_162;
  assign while_if_and_11_cse = NMPRun_wen & while_stage_0_8;
  assign NMP_RunFSM_switch_lp_and_88_cse = NMPRun_wen & and_dcpl_163;
  assign while_if_and_12_cse = NMPRun_wen & while_stage_0_7;
  assign NMP_ComputeSoftmaxExp_for_and_cse = NMPRun_wen & and_dcpl_167 & and_dcpl_164
      & NMP_RunFSM_switch_lp_conc_itm_4_0;
  assign NMP_ComputeSoftmaxExp_for_and_50_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo | reg_max_value_26_0_1_enexo
      | reg_max_value_26_0_enexo | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo |
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo | reg_NMP_ComputeSoftmaxExp_for_asn_30_itm_2_enexo
      | reg_max_value_26_0_sva_dfm_13_1_26_enexo | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo
      | reg_while_stage_0_7_enexo);
  assign NMP_ComputeSoftmaxExp_for_and_51_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_1 | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_1
      | reg_max_value_26_0_enexo_1 | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_1
      | reg_max_value_26_0_1_enexo_1 | reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo
      | reg_max_value_26_0_sva_dfm_13_1_26_enexo_1 | reg_while_stage_0_7_enexo_1
      | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_1);
  assign NMP_ComputeSoftmaxExp_for_and_52_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_max_value_26_0_sva_dfm_13_1_26_enexo_2 | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_2
      | reg_max_value_26_0_1_enexo_2 | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_2
      | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_2 | reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo
      | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_2 | reg_max_value_26_0_enexo_2
      | reg_while_stage_0_7_enexo_2);
  assign NMP_ComputeSoftmaxExp_for_and_53_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_3 | reg_max_value_26_0_enexo_3
      | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_3 | reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo
      | reg_while_stage_0_7_enexo_3 | reg_max_value_26_0_1_enexo_3 | reg_max_value_26_0_sva_dfm_13_1_26_enexo_3
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_3 | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_3);
  assign NMP_ComputeSoftmaxExp_for_and_54_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_while_stage_0_7_enexo_4 | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_4
      | reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo | reg_max_value_26_0_enexo_4
      | reg_max_value_26_0_sva_dfm_13_1_26_enexo_4 | reg_max_value_26_0_1_enexo_4
      | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_4 | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_4
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_4);
  assign NMP_ComputeSoftmaxExp_for_and_55_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_max_value_26_0_enexo_5 | reg_max_value_26_0_sva_dfm_13_1_26_enexo_5
      | reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo | reg_while_stage_0_7_enexo_5
      | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_5 | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_5
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_5 | reg_max_value_26_0_1_enexo_5
      | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_5);
  assign NMP_ComputeSoftmaxExp_for_and_56_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_max_value_26_0_sva_dfm_13_1_26_enexo_6 | reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_2_enexo
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_6 | reg_max_value_26_0_1_enexo_6
      | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_6 | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_6
      | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_6 | reg_max_value_26_0_enexo_6
      | reg_while_stage_0_7_enexo_6);
  assign NMP_ComputeSoftmaxExp_for_and_57_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_2_enexo | reg_max_value_26_0_sva_dfm_13_1_26_enexo_7
      | reg_max_value_26_0_enexo_7 | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_7
      | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_7 | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_7
      | reg_while_stage_0_7_enexo_7 | reg_max_value_26_0_1_enexo_7 | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_7);
  assign NMP_ComputeSoftmaxExp_for_and_58_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_max_value_26_0_1_enexo_8 | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_8
      | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_8 | reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_2_enexo
      | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_8 | reg_max_value_26_0_enexo_8
      | reg_max_value_26_0_sva_dfm_13_1_26_enexo_8 | reg_while_stage_0_7_enexo_8
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_8);
  assign NMP_ComputeSoftmaxExp_for_and_59_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_max_value_26_0_1_enexo_9 | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_9
      | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_9 | reg_max_value_26_0_enexo_9
      | reg_max_value_26_0_sva_dfm_13_1_26_enexo_9 | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_9
      | reg_while_stage_0_7_enexo_9 | reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_2_enexo
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_9);
  assign NMP_ComputeSoftmaxExp_for_and_60_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_max_value_26_0_enexo_10 | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_10
      | reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_2_enexo | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_10
      | reg_while_stage_0_7_enexo_10 | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_10
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_10 | reg_max_value_26_0_1_enexo_10
      | reg_max_value_26_0_sva_dfm_13_1_26_enexo_10);
  assign NMP_ComputeSoftmaxExp_for_and_61_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_11 | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_11
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_11 | reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_2_enexo
      | reg_while_stage_0_7_enexo_11 | reg_max_value_26_0_1_enexo_11 | reg_max_value_26_0_sva_dfm_13_1_26_enexo_11
      | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_11 | reg_max_value_26_0_enexo_11);
  assign NMP_ComputeSoftmaxExp_for_and_62_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_12 | reg_max_value_26_0_sva_dfm_13_1_26_enexo_12
      | reg_while_stage_0_7_enexo_12 | reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_2_enexo
      | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_12 | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_12
      | reg_max_value_26_0_enexo_12 | reg_max_value_26_0_1_enexo_12 | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_12);
  assign NMP_ComputeSoftmaxExp_for_and_63_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_max_value_26_0_1_enexo_13 | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_13
      | reg_max_value_26_0_enexo_13 | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_13
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_13 | reg_while_stage_0_7_enexo_13
      | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_13 | reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_3_enexo
      | reg_max_value_26_0_sva_dfm_13_1_26_enexo_13);
  assign NMP_ComputeSoftmaxExp_for_and_64_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_14 | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_14
      | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_14 | reg_while_stage_0_7_enexo_14
      | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_14 | reg_max_value_26_0_enexo_14
      | reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_3_enexo | reg_max_value_26_0_sva_dfm_13_1_26_enexo_14
      | reg_max_value_26_0_1_enexo_14);
  assign NMP_ComputeSoftmaxExp_for_and_65_enex5 = NMP_ComputeSoftmaxExp_for_and_cse
      & (reg_max_value_26_0_enexo_15 | reg_max_value_26_0_sva_dfm_13_1_26_enexo_15
      | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_15 | reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_15
      | reg_while_stage_0_7_enexo_15 | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_15
      | reg_NMP_ComputeSoftmaxExp_for_asn_itm_3_enexo | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_15
      | reg_max_value_26_0_1_enexo_15);
  assign NMP_RunFSM_switch_lp_and_92_cse = NMPRun_wen & and_dcpl_166;
  assign while_if_and_13_cse = NMPRun_wen & while_stage_0_6;
  assign NMP_RunFSM_switch_lp_and_96_cse = NMPRun_wen & and_dcpl_169;
  assign while_if_and_14_cse = NMPRun_wen & while_stage_0_5;
  assign NMP_RunFSM_switch_lp_and_100_cse = NMPRun_wen & and_dcpl_170;
  assign while_if_and_15_cse = NMPRun_wen & while_stage_0_4;
  assign input_fixed_and_cse = NMPRun_wen & fsm_output;
  assign and_983_cse = input_fixed_and_cse & while_stage_0_4;
  assign NMP_RunFSM_switch_lp_and_104_cse = NMPRun_wen & and_dcpl_171;
  assign input_fixed_and_16_cse = NMPRun_wen & while_stage_0_3;
  assign or_1057_cse = (~(NMP_RunFSM_switch_lp_and_8_cse_1 | NMP_RunFSM_switch_lp_equal_tmp_1))
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign and_1011_cse = (~(or_1057_cse & while_stage_0_4)) & input_fixed_and_16_cse;
  assign and_1236_itm = start_PopNB_mioi_data_rsc_z_mxwt & nmp_config_is_valid_sva;
  assign mux_cse = MUX_s_1_2_2(is_start_sva, and_1236_itm, start_PopNB_mioi_return_rsc_z_mxwt);
  assign nmp_config_num_vector_1_and_cse = NMPRun_wen & (~ or_dcpl_480);
  assign state_and_cse = NMPRun_wen & (~ or_dcpl_481);
  assign nand_7_cse = ~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign while_if_and_17_cse = NMPRun_wen & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign and_1067_cse = (NMP_RunFSM_switch_lp_and_8_cse_1 | NMP_RunFSM_switch_lp_equal_tmp_1)
      & while_stage_0_3 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & NMPRun_wen;
  assign NMP_UpdateFSM_switch_lp_and_4_cse = NMPRun_wen & and_dcpl_172;
  assign large_req_reg_write_data_data_and_112_cse = NMPRun_wen & (~(or_dcpl_679
      | (~ NMP_RunFSM_switch_lp_equal_tmp_9_15) | (~ fsm_output))) & or_dcpl_309;
  assign large_req_reg_write_data_data_and_114_cse = NMPRun_wen & NMP_RunFSM_switch_lp_equal_tmp_9_15
      & (~ or_dcpl_679) & fsm_output & or_dcpl_309;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_cse
      = NMPRun_wen & (~(and_dcpl_634 | or_dcpl_684 | NMP_RunFSM_switch_lp_conc_itm_12_3
      | (~ NMP_RunFSM_switch_lp_conc_itm_12_2) | NMP_RunFSM_switch_lp_conc_itm_12_0));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_5_enex5
      = ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_cse
      & reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_enexo;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_6_enex5
      = ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_cse
      & reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo_2;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_cse
      = NMPRun_wen & (~(((sum_exp_39_4_sva_st_4==36'b000000000000000000000000000000000000))
      | or_dcpl_684 | (~ NMP_RunFSM_switch_lp_conc_itm_12_3) | NMP_RunFSM_switch_lp_conc_itm_12_2
      | NMP_RunFSM_switch_lp_conc_itm_12_0));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5
      = ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_cse
      & reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_5_enex5
      = ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_cse
      & reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_enexo;
  assign nl_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_acc_itm
      = conv_u2u_9_13(ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1[19:11])
      + conv_u2u_12_13({1'b1 , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mux_1_itm_2
      , 1'b1});
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_acc_itm
      = nl_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_acc_itm[12:0];
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_cse = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[33:32]==2'b00)
      & NMP_RunFSM_switch_lp_conc_itm_7_1;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_1_cse = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[33:32]==2'b01)
      & NMP_RunFSM_switch_lp_conc_itm_7_1;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_2_cse = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[33:32]==2'b10)
      & NMP_RunFSM_switch_lp_conc_itm_7_1;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_3_cse = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[33:32]==2'b11)
      & NMP_RunFSM_switch_lp_conc_itm_7_1;
  assign and_1085_enex5 = while_if_and_12_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & (NMP_RunFSM_switch_lp_equal_tmp_5 | NMP_RunFSM_switch_lp_equal_tmp_5_4) &
      (reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_16 | reg_max_value_26_0_sva_dfm_13_1_26_enexo_16
      | reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_16 | reg_max_value_26_0_1_enexo_16
      | reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_16 | reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_16);
  assign NMP_RunFSM_switch_lp_and_126_enex5 = NMPRun_wen & (and_dcpl_292 | and_dcpl_492)
      & reg_NMP_ComputeSoftmaxExp_for_asn_30_itm_2_enexo_1;
  assign max_value_and_1_cse = NMPRun_wen & and_dcpl_292;
  assign NMP_ComputeSoftmaxMax_for_and_enex5 = max_value_and_1_cse & reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo_1;
  assign max_value_and_enex5 = max_value_and_1_cse & (reg_NMP_ComputeSoftmaxMax_for_if_less_5_itm_1_enexo
      | reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo_1 | reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo_1
      | reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo_1 | reg_max_value_26_0_sva_dfm_9_1_26_enexo
      | reg_max_value_26_0_sva_dfm_9_1_25_0_enexo | reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo_1);
  assign NMP_ComputeSoftmaxExp_for_and_66_enex5 = NMP_RunFSM_switch_lp_and_96_cse
      & reg_NMP_RunFSM_switch_lp_asn_104_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_17_cse = NMPRun_wen & (and_dcpl_296 | and_dcpl_342
      | and_dcpl_504);
  assign NMP_ComputeSoftmaxExp_for_and_67_enex5 = NMP_ComputeSoftmaxExp_for_and_17_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_68_enex5 = NMP_ComputeSoftmaxExp_for_and_17_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_69_enex5 = NMP_ComputeSoftmaxExp_for_and_17_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_70_enex5 = NMP_ComputeSoftmaxExp_for_and_17_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_21_enex5 = NMPRun_wen & (and_dcpl_296 | (and_dcpl_346
      & and_dcpl_343 & NMP_ComputeSoftmaxMax_for_if_less_5_tmp) | and_dcpl_504) &
      reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_22_cse = NMPRun_wen & (and_dcpl_296 | and_dcpl_504);
  assign NMP_ComputeSoftmaxExp_for_and_71_enex5 = NMP_ComputeSoftmaxExp_for_and_22_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_72_enex5 = NMP_ComputeSoftmaxExp_for_and_22_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_73_enex5 = NMP_ComputeSoftmaxExp_for_and_22_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_74_enex5 = NMP_ComputeSoftmaxExp_for_and_22_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_75_enex5 = NMP_ComputeSoftmaxExp_for_and_22_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_76_enex5 = NMP_ComputeSoftmaxExp_for_and_22_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_77_enex5 = NMP_ComputeSoftmaxExp_for_and_22_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_29_cse = NMPRun_wen & and_dcpl_296;
  assign NMP_ComputeSoftmaxExp_for_and_78_enex5 = NMP_ComputeSoftmaxExp_for_and_29_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_2_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_79_enex5 = NMP_ComputeSoftmaxExp_for_and_29_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_2_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_80_enex5 = NMP_ComputeSoftmaxExp_for_and_29_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_itm_2_enexo;
  assign or_803_cse = NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign and_899_cse = NMP_RunFSM_switch_lp_or_73_tmp & state_2_sva;
  assign or_801_cse = nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1
      | operator_16_false_acc_2_itm_17;
  assign mux_110_cse = MUX_s_1_2_2(or_tmp_99, mux_tmp_83, or_803_cse);
  assign mux_105_cse_1 = MUX_s_1_2_2(mux_tmp_89, mux_216_itm, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign mux_107_cse = MUX_s_1_2_2(mux_tmp_99, mux_216_itm, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign mux_101_nl = MUX_s_1_2_2(mux_107_cse, mux_105_cse_1, NMP_RunFSM_switch_lp_equal_tmp_11_1);
  assign or_813_nl = (~ NMP_RunFSM_switch_lp_equal_tmp_12_1) | NMP_UpdateFSM_switch_lp_equal_tmp_1
      | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign mux_129_nl = MUX_s_1_2_2(or_tmp_99, mux_tmp_83, or_813_nl);
  assign mux_131_cse = MUX_s_1_2_2(mux_101_nl, mux_129_nl, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_219_cse = MUX_s_1_2_2(mux_tmp_142, nor_tmp_19, or_tmp_129);
  assign mux_216_itm = MUX_s_1_2_2(mux_110_cse, mux_tmp_85, and_899_cse);
  assign or_877_nl = state_3_sva | state_2_sva | not_tmp_279;
  assign or_875_nl = (~ state_3_sva) | state_2_sva | state_0_sva | (~ reg_rva_in_PopNB_mioi_iswt0_cse);
  assign mux_211_nl = MUX_s_1_2_2(or_877_nl, or_875_nl, state_1_sva);
  assign and_896_nl = or_tmp_165 & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign mux_201_nl = MUX_s_1_2_2(and_896_nl, reg_rva_in_PopNB_mioi_iswt0_cse, or_tmp_116);
  assign and_897_nl = next_state_3_lpi_1_dfm_3 & state_2_sva & (~ NMP_RunFSM_switch_lp_equal_tmp_11_1)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign mux_202_nl = MUX_s_1_2_2(mux_201_nl, and_897_nl, NMP_RunFSM_switch_lp_or_73_tmp);
  assign and_673_nl = NMP_RunFSM_switch_lp_equal_tmp_11_1 & not_tmp_286;
  assign mux_199_nl = MUX_s_1_2_2(and_673_nl, reg_rva_in_PopNB_mioi_iswt0_cse, and_899_cse);
  assign mux_203_nl = MUX_s_1_2_2(mux_202_nl, mux_199_nl, state_1_sva_dfm_1);
  assign nand_18_nl = ~(((~(large_rsp_PopNB_mioi_return_rsc_z_mxwt | (~ state_1_sva)))
      | state_3_sva | state_2_sva | state_0_sva) & reg_rva_in_PopNB_mioi_iswt0_cse);
  assign mux_196_nl = MUX_s_1_2_2(nand_18_nl, (~ nor_tmp_31), or_tmp_116);
  assign nor_211_nl = ~(NMP_RunFSM_switch_lp_or_73_tmp | mux_196_nl);
  assign mux_195_nl = MUX_s_1_2_2(not_tmp_286, nor_tmp_31, or_tmp_116);
  assign mux_197_nl = MUX_s_1_2_2(nor_211_nl, mux_195_nl, state_1_sva_dfm_1);
  assign mux_204_nl = MUX_s_1_2_2(mux_203_nl, mux_197_nl, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign nor_212_nl = ~(NMP_RunFSM_switch_lp_equal_tmp_11_1 | or_tmp_159);
  assign mux_191_nl = MUX_s_1_2_2((~ or_tmp_159), nor_212_nl, NMP_RunFSM_switch_lp_or_73_tmp);
  assign mux_192_nl = MUX_s_1_2_2(mux_191_nl, reg_rva_in_PopNB_mioi_iswt0_cse, state_1_sva_dfm_1);
  assign nor_213_nl = ~(NMP_RunFSM_switch_lp_or_73_tmp | nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1
      | operator_16_false_acc_2_itm_17 | not_tmp_279);
  assign or_850_nl = nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1
      | operator_16_false_acc_2_itm_17 | (~ state_1_sva) | (~ state_3_sva) | state_2_sva;
  assign mux_184_nl = MUX_s_1_2_2(not_tmp_277, reg_rva_in_PopNB_mioi_iswt0_cse, or_850_nl);
  assign mux_186_nl = MUX_s_1_2_2(nor_213_nl, mux_184_nl, state_1_sva_dfm_1);
  assign mux_193_nl = MUX_s_1_2_2(mux_192_nl, mux_186_nl, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_205_nl = MUX_s_1_2_2(mux_204_nl, mux_193_nl, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign mux_206_nl = MUX_s_1_2_2(mux_205_nl, (~ or_tmp_147), or_803_cse);
  assign and_901_nl = state_1_sva_dfm_1 & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign mux_207_nl = MUX_s_1_2_2(mux_206_nl, and_901_nl, or_tmp_95);
  assign mux_181_nl = MUX_s_1_2_2((~ or_tmp_147), reg_rva_in_PopNB_mioi_iswt0_cse,
      or_tmp_95);
  assign mux_208_nl = MUX_s_1_2_2(mux_207_nl, mux_181_nl, or_tmp_91);
  assign and_902_nl = or_tmp_92 & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign mux_209_nl = MUX_s_1_2_2(mux_208_nl, and_902_nl, or_tmp_12);
  assign and_903_nl = state_3_sva & state_2_sva;
  assign mux_179_nl = MUX_s_1_2_2(not_tmp_277, reg_rva_in_PopNB_mioi_iswt0_cse, and_903_nl);
  assign and_904_nl = or_tmp & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign mux_180_nl = MUX_s_1_2_2(mux_179_nl, and_904_nl, state_1_sva_dfm_1);
  assign mux_210_nl = MUX_s_1_2_2(mux_209_nl, mux_180_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_212_nl = MUX_s_1_2_2(mux_211_nl, mux_210_nl, while_stage_0_3);
  assign mux_278_nl = MUX_s_1_2_2(mux_110_cse, mux_tmp_85, and_899_cse);
  assign mux_123_nl = MUX_s_1_2_2(mux_278_nl, mux_tmp_85, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign or_811_nl = NMP_RunFSM_switch_lp_equal_tmp_12_1 | NMP_RunFSM_switch_lp_or_73_tmp;
  assign mux_122_nl = MUX_s_1_2_2(mux_110_cse, mux_tmp_85, or_811_nl);
  assign mux_124_nl = MUX_s_1_2_2(mux_123_nl, mux_122_nl, NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2);
  assign mux_126_nl = MUX_s_1_2_2(mux_105_cse_1, mux_124_nl, large_rsp_PopNB_mioi_return_rsc_z_mxwt);
  assign mux_127_nl = MUX_s_1_2_2(mux_107_cse, mux_126_nl, NMP_RunFSM_switch_lp_equal_tmp_11_1);
  assign or_809_nl = (~((~((~ NMP_RunFSM_switch_lp_equal_tmp_11_1) | (~ large_rsp_PopNB_mioi_return_rsc_z_mxwt)
      | NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2)) | NMP_RunFSM_switch_lp_equal_tmp_12_1))
      | NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign mux_121_nl = MUX_s_1_2_2(or_tmp_99, mux_tmp_83, or_809_nl);
  assign mux_128_nl = MUX_s_1_2_2(mux_127_nl, mux_121_nl, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_132_nl = MUX_s_1_2_2(mux_131_cse, mux_128_nl, state_1_sva);
  assign mux_133_nl = MUX_s_1_2_2(mux_132_nl, mux_131_cse, state_0_sva);
  assign mux_134_nl = MUX_s_1_2_2(mux_133_nl, or_tmp_96, or_tmp_95);
  assign mux_115_nl = MUX_s_1_2_2(mux_tmp_99, mux_110_cse, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign mux_112_nl = MUX_s_1_2_2(mux_110_cse, mux_tmp_85, NMP_RunFSM_switch_lp_or_73_tmp);
  assign mux_113_nl = MUX_s_1_2_2(mux_tmp_89, mux_112_nl, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign mux_116_nl = MUX_s_1_2_2(mux_115_nl, mux_113_nl, NMP_RunFSM_switch_lp_equal_tmp_11_1);
  assign mux_117_nl = MUX_s_1_2_2(mux_116_nl, mux_110_cse, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_118_nl = MUX_s_1_2_2(mux_117_nl, mux_131_cse, or_801_cse);
  assign mux_119_nl = MUX_s_1_2_2(mux_131_cse, mux_118_nl, nor_tmp_17);
  assign mux_120_nl = MUX_s_1_2_2(mux_119_nl, or_tmp_96, or_tmp_95);
  assign mux_135_nl = MUX_s_1_2_2(mux_134_nl, mux_120_nl, state_3_sva);
  assign mux_103_nl = MUX_s_1_2_2(mux_131_cse, or_tmp_96, or_tmp_95);
  assign mux_136_nl = MUX_s_1_2_2(mux_135_nl, mux_103_nl, state_2_sva);
  assign or_790_nl = or_tmp_92 | (~ or_tmp_12);
  assign mux_137_nl = MUX_s_1_2_2(mux_136_nl, or_790_nl, or_tmp_91);
  assign mux_81_nl = MUX_s_1_2_2(or_tmp_90, or_tmp_89, state_3_sva);
  assign or_784_nl = state_3_sva | (~ state_0_sva) | state_1_sva_dfm_1;
  assign mux_82_nl = MUX_s_1_2_2(mux_81_nl, or_784_nl, state_2_sva);
  assign mux_138_nl = MUX_s_1_2_2(mux_137_nl, mux_82_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nmp_config_adpbias_1_and_ssc = NMPRun_wen & (~(mux_212_nl & (~((~(mux_138_nl
      & reg_rva_in_PopNB_mioi_iswt0_cse)) & while_stage_0_3))));
  assign and_889_nl = ((~ or_tmp_129) | NMP_UpdateFSM_switch_lp_equal_tmp_4_1 | NMP_UpdateFSM_switch_lp_or_tmp_1)
      & state_1_sva_dfm_1;
  assign mux_149_itm = MUX_s_1_2_2(mux_tmp_147, and_889_nl, next_state_3_lpi_1_dfm_3);
  assign mux_281_nl = MUX_s_1_2_2(mux_tmp_142, nor_tmp_19, or_tmp_129);
  assign mux_146_cse = MUX_s_1_2_2(mux_281_nl, nor_tmp_19, NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2);
  assign sum_exp_and_3_enex5 = NMPRun_wen & and_dcpl_300 & and_dcpl_298 & (~ NMP_RunFSM_switch_lp_conc_itm_8_0)
      & reg_NMP_ComputeSoftmaxSum_for_acc_7_itm_1_enexo;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_6_cse = NMPRun_wen
      & and_dcpl_305 & (~ NMP_RunFSM_switch_lp_conc_itm_6_0) & NMP_RunFSM_switch_lp_conc_itm_6_2
      & (~ NMP_RunFSM_switch_lp_conc_itm_6_3);
  assign NMP_PrepareWriteReq_and_15_cse = NMPRun_wen & and_dcpl_90 & (~ NMP_RunFSM_switch_lp_conc_itm_15_0)
      & NMP_RunFSM_switch_lp_conc_itm_15_1 & NMP_RunFSM_switch_lp_conc_itm_15_3 &
      (~ NMP_RunFSM_switch_lp_conc_itm_15_2);
  assign NMP_ComputeSoftmaxNormalize_for_and_32_cse = NMPRun_wen & and_dcpl_141 &
      and_dcpl_139 & NMP_RunFSM_switch_lp_conc_itm_10_0;
  assign NMP_ComputeSoftmaxNormalize_for_and_96_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_97_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_98_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_99_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_100_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_101_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_102_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_103_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_104_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_105_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_106_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_107_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_108_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_109_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_110_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_111_enex5 = NMP_ComputeSoftmaxNormalize_for_and_32_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_2_enexo;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_2_enex5
      = NMPRun_wen & and_dcpl_317 & (~(NMP_RunFSM_switch_lp_conc_itm_11_1 | NMP_RunFSM_switch_lp_conc_itm_11_2))
      & NMP_RunFSM_switch_lp_conc_itm_11_3 & ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_3
      & NMP_RunFSM_switch_lp_equal_tmp_7_10 & (~ NMP_RunFSM_switch_lp_conc_itm_11_0)
      & reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_enexo;
  assign NMP_ComputeRMSNormalize_for_and_32_cse = NMPRun_wen & and_dcpl_137 & and_dcpl_320;
  assign NMP_ComputeRMSNormalize_for_and_161_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_60_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_162_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_58_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_163_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_56_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_164_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_54_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_165_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_52_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_166_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_50_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_167_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_48_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_168_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_46_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_169_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_44_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_170_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_42_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_171_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_40_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_172_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_38_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_173_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_36_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_174_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_34_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_175_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_32_itm_9_enexo;
  assign NMP_ComputeRMSNormalize_for_and_176_enex5 = NMP_ComputeRMSNormalize_for_and_32_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_itm_9_enexo;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_2_cse = NMPRun_wen
      & and_dcpl_317 & (~ NMP_RunFSM_switch_lp_conc_itm_11_1) & NMP_RunFSM_switch_lp_conc_itm_11_2
      & (~ NMP_RunFSM_switch_lp_conc_itm_11_3) & ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_2_1
      & NMP_RunFSM_switch_lp_equal_tmp_3_10 & (~ NMP_RunFSM_switch_lp_conc_itm_11_0);
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_4_enex5 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_2_cse
      & reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_enexo;
  assign NMP_PrepareReadReq_and_17_cse = NMPRun_wen & and_dcpl_91 & and_dcpl_88 &
      (~ NMP_RunFSM_switch_lp_conc_itm_15_2);
  assign rva_out_reg_data_and_12_cse = NMPRun_wen & while_stage_0_17 & while_while_nor_itm_15;
  assign rva_out_reg_data_and_104_enex5 = rva_out_reg_data_and_12_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_15_enexo;
  assign rva_out_reg_data_and_105_enex5 = rva_out_reg_data_and_12_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_15_enexo;
  assign NMP_RunFSM_switch_lp_and_129_cse = NMPRun_wen & and_dcpl_317;
  assign operator_6_2_true_AC_TRN_AC_WRAP_and_cse = NMPRun_wen & (~(or_dcpl_700 |
      (~(NMP_RunFSM_switch_lp_conc_itm_16_0 & NMP_RunFSM_switch_lp_conc_itm_16_2))
      | NMP_RunFSM_switch_lp_conc_itm_16_3));
  assign operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse = NMPRun_wen & (~(or_dcpl_700
      | (~ NMP_RunFSM_switch_lp_conc_itm_16_0) | NMP_RunFSM_switch_lp_conc_itm_16_2
      | (~ NMP_RunFSM_switch_lp_conc_itm_16_3)));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_1_cse
      = NMPRun_wen & (~(((ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_2==40'b0000000000000000000000000000000000000000))
      | or_dcpl_708 | (~ NMP_RunFSM_switch_lp_conc_itm_11_2) | NMP_RunFSM_switch_lp_conc_itm_11_3
      | NMP_RunFSM_switch_lp_conc_itm_11_0));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_2_cse
      = NMPRun_wen & (~(((sum_exp_39_4_sva_st_3==36'b000000000000000000000000000000000000))
      | or_dcpl_708 | NMP_RunFSM_switch_lp_conc_itm_11_2 | (~ NMP_RunFSM_switch_lp_conc_itm_11_3)
      | NMP_RunFSM_switch_lp_conc_itm_11_0));
  assign sum_exp_and_4_enex5 = NMPRun_wen & ((sum_exp_39_4_sva_st_2!=36'b000000000000000000000000000000000000))
      & and_dcpl_142 & reg_sum_exp_39_4_sva_2_enexo;
  assign NMP_ComputeSoftmaxSum_for_and_cse = NMPRun_wen & and_dcpl_159 & NMP_RunFSM_switch_lp_conc_itm_7_3
      & (~(NMP_RunFSM_switch_lp_conc_itm_7_1 | NMP_RunFSM_switch_lp_conc_itm_7_2
      | NMP_RunFSM_switch_lp_conc_itm_7_0));
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_6_cse
      = NMPRun_wen & ((~ (ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_2[0]))
      | ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_0_3_itm_2)
      & and_dcpl_162 & (~(NMP_RunFSM_switch_lp_conc_itm_6_1 | NMP_RunFSM_switch_lp_conc_itm_6_0))
      & NMP_RunFSM_switch_lp_conc_itm_6_2 & (~ NMP_RunFSM_switch_lp_conc_itm_6_3);
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_8_enex5
      = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_6_cse
      & (reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_enexo
      | reg_NMP_PrepareWriteReq_asn_1_itm_5_1_enexo);
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_9_enex5
      = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_6_cse
      & reg_NMP_PrepareReadReq_asn_2_itm_5_1_enexo;
  assign max_value_and_3_cse = NMPRun_wen & and_dcpl_346 & and_dcpl_343 & (~ NMP_ComputeSoftmaxMax_for_if_less_5_tmp);
  assign max_value_and_9_enex5 = max_value_and_3_cse & (reg_max_value_26_0_sva_dfm_6_1_25_0_enexo
      | reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_1_enexo_1 | reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_1_enexo_1
      | reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_1_enexo_1);
  assign nmp_config_adpbias_1_and_1_ssc = NMPRun_wen & (nmp_config_adpbias_1_sva_dfm_3_1_mx0c0
      | nmp_config_adpbias_1_sva_dfm_3_1_mx0c1 | nmp_config_adpbias_1_sva_dfm_3_1_mx0c2);
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_7_cse = NMPRun_wen
      & and_dcpl_354 & (~(NMP_RunFSM_switch_lp_conc_itm_5_0 | NMP_RunFSM_switch_lp_conc_itm_5_3))
      & NMP_RunFSM_switch_lp_conc_itm_5_2;
  assign NMP_PrepareWriteReq_and_18_cse = NMPRun_wen & and_dcpl_96 & NMP_RunFSM_switch_lp_conc_itm_14_1
      & (~(NMP_RunFSM_switch_lp_conc_itm_14_0 | NMP_RunFSM_switch_lp_conc_itm_14_2))
      & NMP_RunFSM_switch_lp_conc_itm_14_3;
  assign NMP_ComputeSoftmaxNormalize_for_and_48_cse = NMPRun_wen & and_dcpl_365;
  assign NMP_ComputeSoftmaxNormalize_for_and_112_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_113_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_114_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_115_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_116_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_117_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_118_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_119_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_120_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_121_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_122_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_123_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_124_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_125_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_126_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_127_enex5 = NMP_ComputeSoftmaxNormalize_for_and_48_cse
      & reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_32_cse = NMPRun_wen & and_dcpl_367 & (NMP_RunFSM_switch_lp_conc_itm_2_0
      | NMP_RunFSM_switch_lp_conc_itm_2_1) & NMP_RunFSM_switch_lp_conc_itm_2_2;
  assign NMP_ComputeSoftmaxExp_for_and_81_enex5 = NMP_ComputeSoftmaxExp_for_and_32_cse
      & reg_input_fixed_14_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_82_enex5 = NMP_ComputeSoftmaxExp_for_and_32_cse
      & reg_input_fixed_13_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_83_enex5 = NMP_ComputeSoftmaxExp_for_and_32_cse
      & reg_input_fixed_12_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_84_enex5 = NMP_ComputeSoftmaxExp_for_and_32_cse
      & reg_input_fixed_11_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_85_enex5 = NMP_ComputeSoftmaxExp_for_and_32_cse
      & reg_input_fixed_10_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_86_enex5 = NMP_ComputeSoftmaxExp_for_and_32_cse
      & reg_input_fixed_9_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_87_enex5 = NMP_ComputeSoftmaxExp_for_and_32_cse
      & reg_input_fixed_8_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_88_enex5 = NMP_ComputeSoftmaxExp_for_and_32_cse
      & reg_input_fixed_7_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_40_cse = NMPRun_wen & and_dcpl_367 & and_dcpl_369;
  assign NMP_ComputeSoftmaxExp_for_and_89_enex5 = NMP_ComputeSoftmaxExp_for_and_40_cse
      & reg_input_fixed_6_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_90_enex5 = NMP_ComputeSoftmaxExp_for_and_40_cse
      & reg_input_fixed_5_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_91_enex5 = NMP_ComputeSoftmaxExp_for_and_40_cse
      & reg_input_fixed_4_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_92_enex5 = NMP_ComputeSoftmaxExp_for_and_40_cse
      & reg_input_fixed_3_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_44_cse = NMPRun_wen & ((and_dcpl_367 & and_dcpl_369
      & NMP_RunFSM_switch_lp_conc_itm_2_1) | and_dcpl_509);
  assign NMP_ComputeSoftmaxExp_for_and_93_enex5 = NMP_ComputeSoftmaxExp_for_and_44_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_94_enex5 = NMP_ComputeSoftmaxExp_for_and_44_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_1_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_95_enex5 = NMP_ComputeSoftmaxExp_for_and_44_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_itm_1_enexo;
  assign NMP_ComputeRMSNormalize_for_and_48_cse = NMPRun_wen & and_dcpl_377;
  assign NMP_ComputeRMSNormalize_for_and_177_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_60_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_178_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_58_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_179_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_56_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_180_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_54_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_181_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_52_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_182_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_50_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_183_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_48_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_184_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_46_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_185_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_44_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_186_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_42_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_187_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_40_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_188_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_38_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_189_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_36_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_190_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_34_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_191_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_32_itm_8_enexo;
  assign NMP_ComputeRMSNormalize_for_and_192_enex5 = NMP_ComputeRMSNormalize_for_and_48_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_itm_8_enexo;
  assign NMP_PrepareReadReq_and_20_cse = NMPRun_wen & and_dcpl_362 & and_dcpl_360
      & (~ NMP_RunFSM_switch_lp_conc_itm_14_3);
  assign NMP_PrepareReadReq_and_56_enex5 = NMP_PrepareReadReq_and_20_cse & reg_NMP_PrepareReadReq_asn_1_itm_13_1_enexo;
  assign rva_out_reg_data_and_18_cse = NMPRun_wen & while_stage_0_16 & while_while_nor_itm_14;
  assign rva_out_reg_data_and_106_enex5 = rva_out_reg_data_and_18_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_14_enexo;
  assign rva_out_reg_data_and_107_enex5 = rva_out_reg_data_and_18_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_14_enexo;
  assign NMP_RunFSM_switch_lp_and_135_cse = NMPRun_wen & and_dcpl_136 & (~ NMP_RunFSM_switch_lp_equal_tmp_10);
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_13_enex5 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_6_cse
      & reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_2_enexo;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_cse = NMPRun_wen
      & (~(((ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_1==40'b0000000000000000000000000000000000000000))
      | or_dcpl_718 | (~ NMP_RunFSM_switch_lp_conc_itm_10_2) | NMP_RunFSM_switch_lp_conc_itm_10_3
      | NMP_RunFSM_switch_lp_conc_itm_10_1 | NMP_RunFSM_switch_lp_conc_itm_10_0));
  assign nl_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_qif_acc_cse
      = ({1'b1 , (~ rtn_out)}) + 7'b0010001;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_qif_acc_cse = nl_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_qif_acc_cse[6:0];
  assign operator_40_0_false_AC_TRN_AC_WRAP_1_and_enex5 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_cse
      & reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_1_enexo;
  assign sum_exp_and_5_enex5 = NMPRun_wen & reg_sum_exp_39_4_sva_st_1_enexo_1;
  assign and_1094_cse = ((NMP_RunFSM_switch_lp_conc_itm_7_0 & (~ NMP_RunFSM_switch_lp_conc_itm_7_2)
      & (~ NMP_RunFSM_switch_lp_conc_itm_7_1) & NMP_RunFSM_switch_lp_conc_itm_7_3)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | (~ while_stage_0_9) | (~(NMP_RunFSM_switch_lp_equal_tmp_7 | NMP_RunFSM_switch_lp_equal_tmp_6_6)))
      & (NMP_RunFSM_switch_lp_equal_tmp_8 | NMP_RunFSM_switch_lp_equal_tmp_6_7) &
      while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & input_fixed_and_cse;
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_9_cse
      = NMPRun_wen & and_dcpl_159 & NMP_RunFSM_switch_lp_equal_tmp_6_6 & (~ NMP_RunFSM_switch_lp_equal_tmp_7)
      & (~ NMP_RunFSM_switch_lp_conc_itm_7_3) & NMP_RunFSM_switch_lp_conc_itm_7_1
      & NMP_RunFSM_switch_lp_conc_itm_7_2 & NMP_RunFSM_switch_lp_conc_itm_7_0;
  assign and_835_itm = and_dcpl_832 & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_7_cse
      = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[33:32]==2'b00)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_5_cse
      = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[33:32]==2'b10)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_6_cse
      = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[33:32]==2'b11)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign max_value_and_5_cse = NMPRun_wen & and_dcpl_367 & NMP_RunFSM_switch_lp_conc_itm_2_2
      & (~ NMP_RunFSM_switch_lp_conc_itm_2_0) & NMP_RunFSM_switch_lp_conc_itm_2_1;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_9_cse = NMPRun_wen
      & and_dcpl_167 & and_dcpl_409 & (~ NMP_RunFSM_switch_lp_conc_itm_4_0);
  assign NMP_RunFSM_switch_lp_and_342_enex5 = NMP_RunFSM_switch_lp_and_100_cse &
      reg_input_fixed_15_26_0_enexo;
  assign NMP_PrepareWriteReq_and_21_cse = NMPRun_wen & and_dcpl_97 & NMP_RunFSM_switch_lp_conc_itm_13_1
      & (~ NMP_RunFSM_switch_lp_conc_itm_13_0) & NMP_RunFSM_switch_lp_conc_itm_13_3
      & (~ NMP_RunFSM_switch_lp_conc_itm_13_2);
  assign NMP_PrepareWriteReq_and_63_enex5 = NMP_PrepareWriteReq_and_21_cse & reg_NMP_PrepareWriteReq_asn_2_itm_12_enexo;
  assign NMP_PrepareWriteReq_and_64_enex5 = NMP_PrepareWriteReq_and_21_cse & reg_NMP_PrepareWriteReq_asn_2_itm_12_1_enexo;
  assign out_adp_set_value_ac_float_1_and_3_ssc = NMPRun_wen & and_dcpl_418 & NMP_RunFSM_switch_lp_conc_itm_13_0
      & NMP_RunFSM_switch_lp_conc_itm_13_3 & (~ NMP_RunFSM_switch_lp_conc_itm_13_2);
  assign NMP_ComputeSoftmaxNormalize_for_and_64_cse = NMPRun_wen & and_dcpl_300 &
      and_dcpl_298 & NMP_RunFSM_switch_lp_conc_itm_8_0;
  assign NMP_ComputeSoftmaxNormalize_for_and_128_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_15_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_129_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_14_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_130_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_13_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_131_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_12_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_132_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_11_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_133_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_10_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_134_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_9_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_135_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_8_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_136_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_7_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_137_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_6_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_138_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_5_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_139_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_4_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_140_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_3_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_141_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_2_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_142_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_1_enexo;
  assign NMP_ComputeSoftmaxNormalize_for_and_143_enex5 = NMP_ComputeSoftmaxNormalize_for_and_64_cse
      & reg_exp_values_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_47_cse = NMPRun_wen & state_2_sva & state_0_sva
      & (~ state_3_sva) & and_dcpl_171;
  assign NMP_ComputeSoftmaxExp_for_and_96_enex5 = NMP_ComputeSoftmaxExp_for_and_47_cse
      & reg_input_fixed_2_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_97_enex5 = NMP_ComputeSoftmaxExp_for_and_47_cse
      & reg_input_fixed_1_26_0_enexo;
  assign NMP_ComputeSoftmaxExp_for_and_98_enex5 = NMP_ComputeSoftmaxExp_for_and_47_cse
      & reg_input_fixed_0_26_0_enexo;
  assign out_adp_set_value_ac_float_and_3_ssc = NMPRun_wen & and_dcpl_418 & and_dcpl_424
      & NMP_RunFSM_switch_lp_conc_itm_13_2;
  assign NMP_ComputeRMSNormalize_for_and_64_cse = NMPRun_wen & and_dcpl_155 & and_dcpl_427;
  assign NMP_ComputeRMSNormalize_for_and_193_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_60_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_194_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_58_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_195_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_56_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_196_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_54_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_197_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_52_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_198_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_50_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_199_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_48_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_200_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_46_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_201_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_44_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_202_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_42_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_203_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_40_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_204_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_38_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_205_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_36_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_206_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_34_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_207_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_32_itm_7_enexo;
  assign NMP_ComputeRMSNormalize_for_and_208_enex5 = NMP_ComputeRMSNormalize_for_and_64_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_itm_7_enexo;
  assign NMP_PrepareReadReq_and_23_cse = NMPRun_wen & and_dcpl_418 & and_dcpl_424
      & (~ NMP_RunFSM_switch_lp_conc_itm_13_2);
  assign NMP_PrepareReadReq_and_57_enex5 = NMP_PrepareReadReq_and_23_cse & reg_NMP_PrepareReadReq_asn_2_itm_12_1_enexo;
  assign rva_out_reg_data_and_24_cse = NMPRun_wen & while_while_nor_itm_13 & while_stage_0_15;
  assign rva_out_reg_data_and_108_enex5 = rva_out_reg_data_and_24_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_13_enexo;
  assign rva_out_reg_data_and_109_enex5 = rva_out_reg_data_and_24_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_13_enexo;
  assign NMP_RunFSM_switch_lp_and_158_cse = NMPRun_wen & and_dcpl_145 & (~ NMP_RunFSM_switch_lp_equal_tmp_9);
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_14_enex5 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_7_cse
      & reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1_enexo;
  assign nl_NMP_ComputeRMSSqrtRecip_variance_acc_itm = conv_u2u_36_37(sum_sq_1_39_4_sva_mx1)
      + 37'b0000000000000000000000000011010001101;
  assign NMP_ComputeRMSSqrtRecip_variance_acc_itm = nl_NMP_ComputeRMSSqrtRecip_variance_acc_itm[36:0];
  assign max_value_and_7_cse = NMPRun_wen & (~(NMP_ComputeSoftmaxMax_for_if_less_12_tmp
      | state_0_sva)) & state_2_sva & (~ state_3_sva) & and_dcpl_443;
  assign max_value_and_10_enex5 = max_value_and_7_cse & reg_input_fixed_1_26_0_enexo_1;
  assign NMP_PrepareWriteReq_and_24_cse = NMPRun_wen & and_dcpl_100 & NMP_RunFSM_switch_lp_conc_itm_12_1
      & and_dcpl_105 & (~ NMP_RunFSM_switch_lp_conc_itm_12_0);
  assign NMP_ComputeRMSNormalize_for_and_80_cse = NMPRun_wen & and_dcpl_159 & (~
      NMP_RunFSM_switch_lp_conc_itm_7_3) & (~ NMP_RunFSM_switch_lp_conc_itm_7_1)
      & NMP_RunFSM_switch_lp_conc_itm_7_2 & NMP_RunFSM_switch_lp_conc_itm_7_0;
  assign NMP_ComputeRMSNormalize_for_and_209_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_60_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_210_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_58_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_211_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_56_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_212_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_54_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_213_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_52_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_214_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_50_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_215_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_48_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_216_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_46_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_217_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_44_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_218_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_42_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_219_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_40_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_220_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_38_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_221_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_36_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_222_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_34_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_223_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_32_itm_6_enexo;
  assign NMP_ComputeRMSNormalize_for_and_224_enex5 = NMP_ComputeRMSNormalize_for_and_80_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_itm_6_enexo;
  assign NMP_PrepareReadReq_and_26_cse = NMPRun_wen & and_dcpl_101 & (~(NMP_RunFSM_switch_lp_conc_itm_12_3
      | NMP_RunFSM_switch_lp_conc_itm_12_2)) & NMP_RunFSM_switch_lp_conc_itm_12_0;
  assign rva_out_reg_data_and_30_cse = NMPRun_wen & while_while_nor_itm_12 & while_stage_0_14;
  assign rva_out_reg_data_and_110_enex5 = rva_out_reg_data_and_30_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_12_enexo;
  assign rva_out_reg_data_and_111_enex5 = rva_out_reg_data_and_30_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_12_enexo;
  assign NMP_ComputeRMSNormalize_for_and_96_cse = NMPRun_wen & and_dcpl_305 & NMP_RunFSM_switch_lp_conc_itm_6_0
      & NMP_RunFSM_switch_lp_conc_itm_6_2 & (~ NMP_RunFSM_switch_lp_conc_itm_6_3);
  assign NMP_ComputeRMSNormalize_for_and_225_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_60_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_226_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_58_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_227_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_56_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_228_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_54_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_229_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_52_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_230_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_50_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_231_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_48_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_232_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_46_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_233_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_44_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_234_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_42_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_235_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_40_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_236_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_38_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_237_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_36_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_238_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_34_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_239_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_32_itm_5_enexo;
  assign NMP_ComputeRMSNormalize_for_and_240_enex5 = NMP_ComputeRMSNormalize_for_and_96_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_itm_5_enexo;
  assign rva_out_reg_data_and_36_cse = NMPRun_wen & while_while_nor_itm_11 & while_stage_0_13;
  assign rva_out_reg_data_and_112_enex5 = rva_out_reg_data_and_36_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_11_enexo;
  assign rva_out_reg_data_and_113_enex5 = rva_out_reg_data_and_36_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_11_enexo;
  assign NMP_PrepareWriteReq_and_30_ssc = NMPRun_wen & and_dcpl_141 & NMP_RunFSM_switch_lp_conc_itm_10_3
      & NMP_RunFSM_switch_lp_conc_itm_10_1 & (~ NMP_RunFSM_switch_lp_conc_itm_10_0);
  assign NMP_PrepareWriteReq_and_65_enex5 = NMP_PrepareWriteReq_and_30_ssc & reg_NMP_PrepareWriteReq_asn_2_itm_9_enexo;
  assign NMP_PrepareWriteReq_and_66_enex5 = NMP_PrepareWriteReq_and_30_ssc & reg_NMP_PrepareWriteReq_asn_2_itm_9_1_enexo;
  assign NMP_PrepareWriteReq_and_67_enex5 = NMP_PrepareWriteReq_and_30_ssc & reg_NMP_PrepareWriteReq_asn_1_itm_9_2_enexo;
  assign NMP_ComputeRMSNormalize_for_and_112_cse = NMPRun_wen & and_dcpl_354 & and_dcpl_482
      & NMP_RunFSM_switch_lp_conc_itm_5_2;
  assign NMP_ComputeRMSNormalize_for_and_241_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_17;
  assign NMP_ComputeRMSNormalize_for_and_242_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_58_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_243_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_56_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_244_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_54_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_245_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_52_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_246_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_50_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_247_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_48_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_248_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_46_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_249_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_44_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_250_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_42_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_251_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_40_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_252_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_38_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_253_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_36_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_254_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_34_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_255_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_32_itm_4_enexo;
  assign NMP_ComputeRMSNormalize_for_and_256_enex5 = NMP_ComputeRMSNormalize_for_and_112_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_itm_4_enexo;
  assign NMP_PrepareReadReq_and_32_ssc = NMPRun_wen & and_dcpl_141 & and_dcpl_320;
  assign NMP_PrepareReadReq_and_58_enex5 = NMP_PrepareReadReq_and_32_ssc & reg_NMP_PrepareReadReq_asn_2_itm_9_enexo;
  assign NMP_PrepareReadReq_and_59_enex5 = NMP_PrepareReadReq_and_32_ssc & reg_NMP_PrepareReadReq_asn_2_itm_9_1_enexo;
  assign xor_3_ssc = NMP_RunFSM_switch_lp_conc_itm_10_2 ^ NMP_RunFSM_switch_lp_conc_itm_10_3;
  assign rva_out_reg_data_and_42_cse = NMPRun_wen & while_stage_0_12 & while_while_nor_itm_10;
  assign rva_out_reg_data_and_114_enex5 = rva_out_reg_data_and_42_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_10_enexo;
  assign rva_out_reg_data_and_115_enex5 = rva_out_reg_data_and_42_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_10_enexo;
  assign NMP_PrepareWriteReq_and_35_cse = NMPRun_wen & and_dcpl_150 & NMP_RunFSM_switch_lp_conc_itm_9_3
      & NMP_RunFSM_switch_lp_conc_itm_9_1 & (~ NMP_RunFSM_switch_lp_conc_itm_9_0);
  assign NMP_ComputeRMSNormalize_for_and_128_cse = NMPRun_wen & and_dcpl_492;
  assign NMP_ComputeRMSNormalize_for_and_257_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo_2;
  assign NMP_ComputeRMSNormalize_for_and_258_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo_2;
  assign NMP_ComputeRMSNormalize_for_and_259_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo_2;
  assign NMP_ComputeRMSNormalize_for_and_260_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo_2;
  assign NMP_ComputeRMSNormalize_for_and_261_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo_2;
  assign NMP_ComputeRMSNormalize_for_and_262_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_2_enexo_1;
  assign NMP_ComputeRMSNormalize_for_and_263_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_2_enexo_1;
  assign NMP_ComputeRMSNormalize_for_and_264_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_2_enexo_1;
  assign NMP_ComputeRMSNormalize_for_and_265_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_2_enexo_1;
  assign NMP_ComputeRMSNormalize_for_and_266_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_2_enexo_1;
  assign NMP_ComputeRMSNormalize_for_and_267_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_2_enexo_1;
  assign NMP_ComputeRMSNormalize_for_and_268_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_2_enexo_1;
  assign NMP_ComputeRMSNormalize_for_and_269_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_34_itm_3_enexo;
  assign NMP_ComputeRMSNormalize_for_and_270_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_1_enexo;
  assign NMP_ComputeRMSNormalize_for_and_271_enex5 = NMP_ComputeRMSNormalize_for_and_128_cse
      & reg_NMP_ComputeRMSNormalize_for_asn_itm_3_enexo;
  assign NMP_PrepareReadReq_and_36_cse = NMPRun_wen & and_dcpl_150 & and_dcpl_376;
  assign rva_out_reg_data_and_48_cse = NMPRun_wen & while_stage_0_11 & while_while_nor_itm_9;
  assign rva_out_reg_data_and_116_enex5 = rva_out_reg_data_and_48_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_9_enexo;
  assign rva_out_reg_data_and_117_enex5 = rva_out_reg_data_and_48_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_9_enexo;
  assign NMP_PrepareWriteReq_and_38_cse = NMPRun_wen & and_dcpl_300 & NMP_RunFSM_switch_lp_conc_itm_8_1
      & NMP_RunFSM_switch_lp_conc_itm_8_3 & (~ NMP_RunFSM_switch_lp_conc_itm_8_0);
  assign NMP_ComputeRMSNormalize_for_and_143_cse = NMPRun_wen & and_dcpl_504;
  assign NMP_ComputeRMSNormalize_for_and_272_enex5 = NMP_ComputeRMSNormalize_for_and_143_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_2_enexo_1;
  assign NMP_ComputeRMSNormalize_for_and_273_enex5 = NMP_ComputeRMSNormalize_for_and_143_cse
      & reg_NMP_ComputeSoftmaxExp_for_asn_itm_2_enexo_1;
  assign NMP_PrepareReadReq_and_39_cse = NMPRun_wen & and_dcpl_300 & and_dcpl_427;
  assign rva_out_reg_data_and_54_cse = NMPRun_wen & while_stage_0_10 & while_while_nor_itm_8;
  assign rva_out_reg_data_and_118_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_8_enexo;
  assign rva_out_reg_data_and_119_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_8_enexo;
  assign rva_out_reg_data_and_60_cse = NMPRun_wen & while_while_nor_itm_7 & while_stage_0_9;
  assign rva_out_reg_data_and_120_enex5 = rva_out_reg_data_and_60_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_7_enexo;
  assign rva_out_reg_data_and_121_enex5 = rva_out_reg_data_and_60_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_7_enexo;
  assign NMP_PrepareWriteReq_and_41_cse = NMPRun_wen & and_dcpl_162 & NMP_RunFSM_switch_lp_conc_itm_6_1
      & (~(NMP_RunFSM_switch_lp_conc_itm_6_0 | NMP_RunFSM_switch_lp_conc_itm_6_2))
      & NMP_RunFSM_switch_lp_conc_itm_6_3;
  assign NMP_PrepareWriteReq_and_68_enex5 = NMP_PrepareWriteReq_and_41_cse & reg_NMP_PrepareWriteReq_asn_2_itm_5_enexo;
  assign NMP_PrepareReadReq_and_44_cse = NMPRun_wen & and_dcpl_305 & and_dcpl_519
      & (~ NMP_RunFSM_switch_lp_conc_itm_6_3);
  assign rva_out_reg_data_and_66_cse = NMPRun_wen & while_while_nor_itm_6 & while_stage_0_8;
  assign rva_out_reg_data_and_122_enex5 = rva_out_reg_data_and_66_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_6_enexo;
  assign rva_out_reg_data_and_123_enex5 = rva_out_reg_data_and_66_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_6_enexo;
  assign NMP_PrepareWriteReq_and_44_cse = NMPRun_wen & and_dcpl_163 & NMP_RunFSM_switch_lp_conc_itm_5_1
      & (~ NMP_RunFSM_switch_lp_conc_itm_5_0) & NMP_RunFSM_switch_lp_conc_itm_5_3
      & (~ NMP_RunFSM_switch_lp_conc_itm_5_2);
  assign NMP_PrepareWriteReq_and_69_enex5 = NMP_PrepareWriteReq_and_44_cse & reg_NMP_PrepareWriteReq_asn_2_itm_4_enexo;
  assign NMP_PrepareWriteReq_and_8_cse = (operator_40_0_false_AC_TRN_AC_WRAP_lshift_itm[38:37]==2'b00)
      & NMP_RunFSM_switch_lp_conc_itm_5_2;
  assign NMP_PrepareWriteReq_and_9_cse = (operator_40_0_false_AC_TRN_AC_WRAP_lshift_itm[38:37]==2'b01)
      & NMP_RunFSM_switch_lp_conc_itm_5_2;
  assign NMP_PrepareWriteReq_and_10_cse = (operator_40_0_false_AC_TRN_AC_WRAP_lshift_itm[38:37]==2'b10)
      & NMP_RunFSM_switch_lp_conc_itm_5_2;
  assign NMP_PrepareWriteReq_and_11_cse = (operator_40_0_false_AC_TRN_AC_WRAP_lshift_itm[38:37]==2'b11)
      & NMP_RunFSM_switch_lp_conc_itm_5_2;
  assign rva_out_reg_data_and_72_cse = NMPRun_wen & while_stage_0_7 & while_while_nor_itm_5;
  assign rva_out_reg_data_and_124_enex5 = rva_out_reg_data_and_72_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_5_enexo;
  assign rva_out_reg_data_and_125_enex5 = rva_out_reg_data_and_72_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_5_enexo;
  assign NMP_PrepareWriteReq_and_47_cse = NMPRun_wen & and_dcpl_541 & (~ NMP_RunFSM_switch_lp_conc_itm_4_2)
      & NMP_RunFSM_switch_lp_conc_itm_4_1 & (~ NMP_RunFSM_switch_lp_conc_itm_4_0);
  assign NMP_PrepareWriteReq_and_70_enex5 = NMP_PrepareWriteReq_and_47_cse & reg_NMP_PrepareWriteReq_asn_2_itm_3_enexo;
  assign NMP_PrepareWriteReq_and_71_enex5 = NMP_PrepareWriteReq_and_47_cse & reg_NMP_PrepareWriteReq_asn_1_itm_3_enexo;
  assign out_adp_set_value_ac_float_1_and_11_ssc = NMPRun_wen & and_dcpl_541 & and_dcpl_544;
  assign NMP_PrepareReadReq_and_47_cse = NMPRun_wen & and_dcpl_167 & and_dcpl_544;
  assign NMP_PrepareReadReq_and_60_enex5 = NMP_PrepareReadReq_and_47_cse & reg_NMP_PrepareReadReq_asn_2_itm_3_enexo;
  assign rva_out_reg_data_and_78_cse = NMPRun_wen & while_while_nor_itm_4 & while_stage_0_6;
  assign rva_out_reg_data_and_126_enex5 = rva_out_reg_data_and_78_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_4_enexo;
  assign rva_out_reg_data_and_127_enex5 = rva_out_reg_data_and_78_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_4_enexo;
  assign NMP_PrepareWriteReq_and_50_cse = NMPRun_wen & and_dcpl_554 & (~ NMP_RunFSM_switch_lp_conc_itm_3_2)
      & NMP_RunFSM_switch_lp_conc_itm_3_1 & (~ NMP_RunFSM_switch_lp_conc_itm_3_0);
  assign NMP_PrepareWriteReq_and_72_enex5 = NMP_PrepareWriteReq_and_50_cse & reg_NMP_PrepareWriteReq_asn_2_itm_2_enexo;
  assign NMP_PrepareWriteReq_and_73_enex5 = NMP_PrepareWriteReq_and_50_cse & reg_NMP_PrepareWriteReq_asn_1_itm_2_enexo;
  assign NMP_PrepareReadReq_and_50_cse = NMPRun_wen & and_dcpl_295 & and_dcpl_557;
  assign NMP_PrepareReadReq_and_61_enex5 = NMP_PrepareReadReq_and_50_cse & reg_NMP_PrepareWriteReq_asn_2_itm_2_enexo_1;
  assign NMP_PrepareReadReq_and_62_enex5 = NMP_PrepareReadReq_and_50_cse & reg_NMP_PrepareWriteReq_asn_1_itm_2_enexo_1;
  assign rva_out_reg_data_and_84_cse = NMPRun_wen & while_while_nor_itm_3 & while_stage_0_5;
  assign rva_out_reg_data_and_128_enex5 = rva_out_reg_data_and_84_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_3_enexo;
  assign rva_out_reg_data_and_129_enex5 = rva_out_reg_data_and_84_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_3_enexo;
  assign NMP_PrepareWriteReq_and_53_cse = NMPRun_wen & ((and_dcpl_564 & (~(NMP_RunFSM_switch_lp_conc_itm_2_2
      | NMP_RunFSM_switch_lp_conc_itm_2_0)) & NMP_RunFSM_switch_lp_conc_itm_2_1)
      | (and_dcpl_367 & and_dcpl_567));
  assign NMP_PrepareWriteReq_and_74_enex5 = NMP_PrepareWriteReq_and_53_cse & reg_NMP_PrepareWriteReq_asn_2_itm_1_enexo;
  assign NMP_PrepareWriteReq_and_75_enex5 = NMP_PrepareWriteReq_and_53_cse & reg_NMP_PrepareWriteReq_asn_1_itm_1_enexo;
  assign rva_out_reg_data_and_90_cse = NMPRun_wen & while_stage_0_4 & while_while_nor_itm_2;
  assign rva_out_reg_data_and_130_enex5 = rva_out_reg_data_and_90_cse & reg_rva_out_reg_data_79_64_sva_dfm_3_2_enexo;
  assign rva_out_reg_data_and_131_enex5 = rva_out_reg_data_and_90_cse & reg_rva_out_reg_data_55_48_sva_dfm_3_2_enexo;
  assign nor_66_nl = ~(state_3_sva | (~ state_0_sva));
  assign nor_67_nl = ~((~ state_3_sva) | state_0_sva);
  assign mux_15_nl = MUX_s_1_2_2(nor_66_nl, nor_67_nl, state_1_sva);
  assign NMP_PrepareWriteReq_and_56_cse = NMPRun_wen & mux_15_nl & (~(state_2_sva
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign NMP_PrepareWriteReq_and_76_enex5 = NMP_PrepareWriteReq_and_56_cse & reg_nmp_config_timestep_counter_enexo;
  assign NMP_PrepareWriteReq_and_77_enex5 = NMP_PrepareWriteReq_and_56_cse & reg_nmp_config_vector_counter_enexo;
  assign rva_out_reg_data_and_96_cse = NMPRun_wen & while_while_nor_itm_1 & while_stage_0_3;
  assign rva_out_reg_data_and_132_enex5 = rva_out_reg_data_and_96_cse & reg_rva_out_reg_data_79_64_enexo;
  assign rva_out_reg_data_and_133_enex5 = rva_out_reg_data_and_96_cse & reg_rva_out_reg_data_55_48_enexo;
  assign or_503_cse = (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign while_and_142_rgt = and_dcpl_875 & (~ or_503_cse);
  assign rva_out_reg_data_and_1_cse = NMPRun_wen & and_dcpl_875 & (~(nand_7_cse |
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
  assign input_fixed_mux_1_cse = MUX_v_27_2_2(input_fixed_12_26_0_sva, input_fixed_12_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_3_cse = MUX_v_27_2_2(input_fixed_13_26_0_sva, input_fixed_13_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_5_cse = MUX_v_27_2_2(input_fixed_14_26_0_sva, input_fixed_14_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_7_cse = MUX_v_27_2_2(input_fixed_15_26_0_sva, input_fixed_15_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_9_cse = MUX_v_27_2_2(input_fixed_3_26_0_sva, input_fixed_3_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_11_cse = MUX_v_27_2_2(input_fixed_4_26_0_sva, input_fixed_4_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_13_cse = MUX_v_27_2_2(input_fixed_5_26_0_sva, input_fixed_5_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_15_cse = MUX_v_27_2_2(input_fixed_6_26_0_sva, input_fixed_6_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_17_cse = MUX_v_27_2_2(input_fixed_7_26_0_sva, input_fixed_7_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_19_cse = MUX_v_27_2_2(input_fixed_8_26_0_sva, input_fixed_8_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_21_cse = MUX_v_27_2_2(input_fixed_9_26_0_sva, input_fixed_9_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_23_cse = MUX_v_27_2_2(input_fixed_10_26_0_sva, input_fixed_10_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign input_fixed_mux_25_cse = MUX_v_27_2_2(input_fixed_11_26_0_sva, input_fixed_11_26_0_sva_dfm_2_1,
      while_stage_0_4);
  assign write_data_data_15_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_15_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_15_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_15_3_0_sva_dfm_1,
      write_data_data_15_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_14_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_14_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_15_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_15_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_14_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_14_3_0_sva_dfm_1,
      write_data_data_14_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_13_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_13_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_14_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_14_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_13_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_13_3_0_sva_dfm_1,
      write_data_data_13_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_12_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_12_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_13_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_13_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_12_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_12_3_0_sva_dfm_1,
      write_data_data_12_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_11_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_11_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_12_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_12_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_11_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_11_3_0_sva_dfm_1,
      write_data_data_11_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_10_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_10_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_11_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_11_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_10_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_10_3_0_sva_dfm_1,
      write_data_data_10_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_9_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_9_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_10_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_10_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_9_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_9_3_0_sva_dfm_1,
      write_data_data_9_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_8_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_8_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_9_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_9_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_8_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_8_3_0_sva_dfm_1,
      write_data_data_8_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_7_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_7_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_8_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_8_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_7_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_7_3_0_sva_dfm_1,
      write_data_data_7_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_6_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_6_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_7_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_7_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_6_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_6_3_0_sva_dfm_1,
      write_data_data_6_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_5_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_5_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_6_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_6_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_5_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_5_3_0_sva_dfm_1,
      write_data_data_5_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_4_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_4_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_5_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_5_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_4_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_4_3_0_sva_dfm_1,
      write_data_data_4_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_3_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_3_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_4_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_4_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_3_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_3_3_0_sva_dfm_1,
      write_data_data_3_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_2_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_2_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_3_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_3_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_2_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_2_3_0_sva_dfm_1,
      write_data_data_2_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_1_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_1_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_2_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_2_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_1_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_1_3_0_sva_dfm_1,
      write_data_data_1_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign write_data_data_0_3_0_sva_dfm_1_mx0w0 = MUX1HOT_v_4_3_2(write_data_data_0_3_0_sva_dfm_1,
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_1_lpi_1_dfm_1_1, NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_1_lpi_1_dfm_1_1,
      {while_asn_728 , while_asn_730 , while_asn_732});
  assign write_data_data_0_3_0_sva_dfm_1_mx1 = MUX_v_4_2_2(write_data_data_0_3_0_sva_dfm_1,
      write_data_data_0_3_0_sva_dfm_1_mx0w0, while_stage_0_20);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_45_nl = out_float_round_32_if_m_1_1_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_45_nl = out_float_round_32_1_if_m_1_1_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_905_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_15_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_45_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_45_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign operator_5_true_not_110_nl = ~ NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_32_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_110_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_32_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_32_nl, 2'b11, out_adp_set_value_ac_float_lor_lpi_1_dfm_1));
  assign operator_5_true_1_not_110_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_32_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_110_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_32_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_32_nl, 2'b11, out_adp_set_value_ac_float_1_lor_lpi_1_dfm_1));
  assign write_data_data_15_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_15_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_32_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_32_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_75_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_668_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_16_itm_1
      | out_adp_set_value_ac_float_mux_95_tmp_3;
  assign operator_5_true_mux_31_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_668_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_15_nl
      = ~((~(out_adp_set_value_ac_float_mux_75_nl | (~ operator_5_true_mux_31_nl)))
      | out_adp_set_value_ac_float_lor_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_75_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_766_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_16_itm_1
      | out_adp_set_value_ac_float_1_mux_95_tmp_3;
  assign operator_5_true_1_mux_31_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_766_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_15_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_75_nl | (~ operator_5_true_1_mux_31_nl)))
      | out_adp_set_value_ac_float_1_lor_lpi_1_dfm_1);
  assign write_data_data_15_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_15_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_15_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_15_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign operator_5_true_not_80_nl = ~ NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_33_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_1_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_80_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_33_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_33_nl, 2'b11, out_adp_set_value_ac_float_lor_1_lpi_1_dfm_1));
  assign operator_5_true_1_not_80_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_33_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_1_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_80_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_33_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_33_nl, 2'b11, out_adp_set_value_ac_float_1_lor_1_lpi_1_dfm_1));
  assign write_data_data_0_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_0_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_33_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_33_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_1_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_1_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_578_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_itm_1
      | out_adp_set_value_ac_float_mux_80_tmp_3;
  assign operator_5_true_mux_1_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_578_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_nl
      = ~((~(out_adp_set_value_ac_float_mux_nl | (~ operator_5_true_mux_1_nl))) |
      out_adp_set_value_ac_float_lor_1_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_1_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_1_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_676_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1
      | out_adp_set_value_ac_float_1_mux_80_tmp_3;
  assign operator_5_true_1_mux_1_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_676_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_nl | (~ operator_5_true_1_mux_1_nl)))
      | out_adp_set_value_ac_float_1_lor_1_lpi_1_dfm_1);
  assign write_data_data_0_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_0_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_nl = out_float_round_32_if_m_1_3_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_1_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_nl = out_float_round_32_1_if_m_1_3_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_1_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_860_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_0_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_42_nl = out_float_round_32_if_m_1_17_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_15_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_42_nl = out_float_round_32_1_if_m_1_17_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_15_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_902_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_14_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_42_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_42_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign operator_5_true_not_108_nl = ~ NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_34_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_15_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_108_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_34_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_34_nl, 2'b11, out_adp_set_value_ac_float_lor_15_lpi_1_dfm_1));
  assign operator_5_true_1_not_108_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_34_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_15_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_108_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_34_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_34_nl, 2'b11, out_adp_set_value_ac_float_1_lor_15_lpi_1_dfm_1));
  assign write_data_data_14_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_14_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_34_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_34_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_70_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_15_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_15_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_662_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1
      | out_adp_set_value_ac_float_mux_94_tmp_3;
  assign operator_5_true_mux_29_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_662_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_14_nl
      = ~((~(out_adp_set_value_ac_float_mux_70_nl | (~ operator_5_true_mux_29_nl)))
      | out_adp_set_value_ac_float_lor_15_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_70_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_15_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_15_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_760_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_15_itm_1
      | out_adp_set_value_ac_float_1_mux_94_tmp_3;
  assign operator_5_true_1_mux_29_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_760_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_14_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_70_nl | (~ operator_5_true_1_mux_29_nl)))
      | out_adp_set_value_ac_float_1_lor_15_lpi_1_dfm_1);
  assign write_data_data_14_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_14_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_14_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_14_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign operator_5_true_not_82_nl = ~ NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_35_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_2_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_82_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_35_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_35_nl, 2'b11, out_adp_set_value_ac_float_lor_2_lpi_1_dfm_1));
  assign operator_5_true_1_not_82_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_35_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_2_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_82_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_35_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_35_nl, 2'b11, out_adp_set_value_ac_float_1_lor_2_lpi_1_dfm_1));
  assign write_data_data_1_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_1_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_35_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_35_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_5_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_2_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_2_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_584_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_2_itm_1
      | out_adp_set_value_ac_float_mux_81_tmp_3;
  assign operator_5_true_mux_3_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_584_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_1_nl
      = ~((~(out_adp_set_value_ac_float_mux_5_nl | (~ operator_5_true_mux_3_nl)))
      | out_adp_set_value_ac_float_lor_2_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_5_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_2_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_2_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_682_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1
      | out_adp_set_value_ac_float_1_mux_81_tmp_3;
  assign operator_5_true_1_mux_3_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_682_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_1_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_5_nl | (~ operator_5_true_1_mux_3_nl)))
      | out_adp_set_value_ac_float_1_lor_2_lpi_1_dfm_1);
  assign write_data_data_1_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_1_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_1_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_1_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_3_nl = out_float_round_32_if_m_1_4_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_2_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_3_nl = out_float_round_32_1_if_m_1_4_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_2_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_863_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_1_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_3_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_3_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_39_nl = out_float_round_32_if_m_1_16_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_14_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_39_nl = out_float_round_32_1_if_m_1_16_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_14_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_899_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_13_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_39_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_39_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign operator_5_true_not_106_nl = ~ NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_36_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_14_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_106_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_36_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_36_nl, 2'b11, out_adp_set_value_ac_float_lor_14_lpi_1_dfm_1));
  assign operator_5_true_1_not_106_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_36_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_14_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_106_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_36_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_36_nl, 2'b11, out_adp_set_value_ac_float_1_lor_14_lpi_1_dfm_1));
  assign write_data_data_13_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_13_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_36_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_36_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_65_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_14_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_14_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_656_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_14_itm_1
      | out_adp_set_value_ac_float_mux_93_tmp_3;
  assign operator_5_true_mux_27_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_656_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_13_nl
      = ~((~(out_adp_set_value_ac_float_mux_65_nl | (~ operator_5_true_mux_27_nl)))
      | out_adp_set_value_ac_float_lor_14_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_65_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_14_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_14_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_754_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1
      | out_adp_set_value_ac_float_1_mux_93_tmp_3;
  assign operator_5_true_1_mux_27_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_754_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_13_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_65_nl | (~ operator_5_true_1_mux_27_nl)))
      | out_adp_set_value_ac_float_1_lor_14_lpi_1_dfm_1);
  assign write_data_data_13_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_13_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_13_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_13_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign operator_5_true_not_84_nl = ~ NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_37_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_3_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_84_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_37_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_37_nl, 2'b11, out_adp_set_value_ac_float_lor_3_lpi_1_dfm_1));
  assign operator_5_true_1_not_84_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_37_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_3_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_84_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_37_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_37_nl, 2'b11, out_adp_set_value_ac_float_1_lor_3_lpi_1_dfm_1));
  assign write_data_data_2_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_2_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_37_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_37_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_10_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_3_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_3_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_590_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_3_itm_1
      | out_adp_set_value_ac_float_mux_82_tmp_3;
  assign operator_5_true_mux_5_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_590_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_2_nl
      = ~((~(out_adp_set_value_ac_float_mux_10_nl | (~ operator_5_true_mux_5_nl)))
      | out_adp_set_value_ac_float_lor_3_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_10_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_3_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_3_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_688_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1
      | out_adp_set_value_ac_float_1_mux_82_tmp_3;
  assign operator_5_true_1_mux_5_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_688_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_2_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_10_nl | (~ operator_5_true_1_mux_5_nl)))
      | out_adp_set_value_ac_float_1_lor_3_lpi_1_dfm_1);
  assign write_data_data_2_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_2_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_2_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_2_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_6_nl = out_float_round_32_if_m_1_5_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_3_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_6_nl = out_float_round_32_1_if_m_1_5_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_3_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_866_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_2_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_6_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_6_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_36_nl = out_float_round_32_if_m_1_15_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_13_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_36_nl = out_float_round_32_1_if_m_1_15_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_13_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_896_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_12_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_36_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_36_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign operator_5_true_not_104_nl = ~ NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_38_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_13_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_104_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_38_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_38_nl, 2'b11, out_adp_set_value_ac_float_lor_13_lpi_1_dfm_1));
  assign operator_5_true_1_not_104_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_38_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_13_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_104_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_38_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_38_nl, 2'b11, out_adp_set_value_ac_float_1_lor_13_lpi_1_dfm_1));
  assign write_data_data_12_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_12_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_38_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_38_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_60_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_13_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_13_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_650_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_13_itm_1
      | out_adp_set_value_ac_float_mux_92_tmp_3;
  assign operator_5_true_mux_25_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_650_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_12_nl
      = ~((~(out_adp_set_value_ac_float_mux_60_nl | (~ operator_5_true_mux_25_nl)))
      | out_adp_set_value_ac_float_lor_13_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_60_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_13_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_13_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_748_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_13_itm_1
      | out_adp_set_value_ac_float_1_mux_92_tmp_3;
  assign operator_5_true_1_mux_25_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_748_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_12_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_60_nl | (~ operator_5_true_1_mux_25_nl)))
      | out_adp_set_value_ac_float_1_lor_13_lpi_1_dfm_1);
  assign write_data_data_12_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_12_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_12_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_12_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign operator_5_true_not_86_nl = ~ NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_39_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_4_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_86_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_39_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_39_nl, 2'b11, out_adp_set_value_ac_float_lor_4_lpi_1_dfm_1));
  assign operator_5_true_1_not_86_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_39_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_4_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_86_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_39_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_39_nl, 2'b11, out_adp_set_value_ac_float_1_lor_4_lpi_1_dfm_1));
  assign write_data_data_3_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_3_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_39_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_39_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_15_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_4_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_4_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_596_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_4_itm_1
      | out_adp_set_value_ac_float_mux_83_tmp_3;
  assign operator_5_true_mux_7_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_596_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_3_nl
      = ~((~(out_adp_set_value_ac_float_mux_15_nl | (~ operator_5_true_mux_7_nl)))
      | out_adp_set_value_ac_float_lor_4_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_15_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_4_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_4_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_694_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1
      | out_adp_set_value_ac_float_1_mux_83_tmp_3;
  assign operator_5_true_1_mux_7_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_694_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_3_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_15_nl | (~ operator_5_true_1_mux_7_nl)))
      | out_adp_set_value_ac_float_1_lor_4_lpi_1_dfm_1);
  assign write_data_data_3_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_3_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_3_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_3_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_9_nl = out_float_round_32_if_m_1_6_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_4_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_9_nl = out_float_round_32_1_if_m_1_6_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_4_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_869_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_3_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_9_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_9_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_33_nl = out_float_round_32_if_m_1_14_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_12_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_33_nl = out_float_round_32_1_if_m_1_14_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_12_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_893_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_11_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_33_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_33_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign operator_5_true_not_102_nl = ~ NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_40_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_12_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_102_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_40_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_40_nl, 2'b11, out_adp_set_value_ac_float_lor_12_lpi_1_dfm_1));
  assign operator_5_true_1_not_102_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_40_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_12_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_102_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_40_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_40_nl, 2'b11, out_adp_set_value_ac_float_1_lor_12_lpi_1_dfm_1));
  assign write_data_data_11_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_11_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_40_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_40_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_55_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_12_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_12_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_644_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1
      | out_adp_set_value_ac_float_mux_91_tmp_3;
  assign operator_5_true_mux_23_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_644_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_11_nl
      = ~((~(out_adp_set_value_ac_float_mux_55_nl | (~ operator_5_true_mux_23_nl)))
      | out_adp_set_value_ac_float_lor_12_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_55_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_12_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_12_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_742_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_12_itm_1
      | out_adp_set_value_ac_float_1_mux_91_tmp_3;
  assign operator_5_true_1_mux_23_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_742_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_11_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_55_nl | (~ operator_5_true_1_mux_23_nl)))
      | out_adp_set_value_ac_float_1_lor_12_lpi_1_dfm_1);
  assign write_data_data_11_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_11_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_11_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_11_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign operator_5_true_not_88_nl = ~ NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_41_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_5_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_88_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_41_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_41_nl, 2'b11, out_adp_set_value_ac_float_lor_5_lpi_1_dfm_1));
  assign operator_5_true_1_not_88_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_41_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_5_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_88_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_41_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_41_nl, 2'b11, out_adp_set_value_ac_float_1_lor_5_lpi_1_dfm_1));
  assign write_data_data_4_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_4_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_41_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_41_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_20_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_5_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_5_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_602_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1
      | out_adp_set_value_ac_float_mux_84_tmp_3;
  assign operator_5_true_mux_9_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_602_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_4_nl
      = ~((~(out_adp_set_value_ac_float_mux_20_nl | (~ operator_5_true_mux_9_nl)))
      | out_adp_set_value_ac_float_lor_5_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_20_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_5_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_5_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_700_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_5_itm_1
      | out_adp_set_value_ac_float_1_mux_84_tmp_3;
  assign operator_5_true_1_mux_9_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_700_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_4_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_20_nl | (~ operator_5_true_1_mux_9_nl)))
      | out_adp_set_value_ac_float_1_lor_5_lpi_1_dfm_1);
  assign write_data_data_4_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_4_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_4_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_4_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_12_nl = out_float_round_32_if_m_1_7_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_5_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_12_nl = out_float_round_32_1_if_m_1_7_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_5_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_872_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_4_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_12_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_12_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_30_nl = out_float_round_32_if_m_1_13_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_11_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_30_nl = out_float_round_32_1_if_m_1_13_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_11_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_890_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_10_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_30_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_30_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign operator_5_true_not_100_nl = ~ NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_42_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_11_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_100_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_42_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_42_nl, 2'b11, out_adp_set_value_ac_float_lor_11_lpi_1_dfm_1));
  assign operator_5_true_1_not_100_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_42_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_11_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_100_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_42_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_42_nl, 2'b11, out_adp_set_value_ac_float_1_lor_11_lpi_1_dfm_1));
  assign write_data_data_10_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_10_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_42_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_42_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_50_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_11_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_11_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_638_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1
      | out_adp_set_value_ac_float_mux_90_tmp_3;
  assign operator_5_true_mux_21_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_638_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_10_nl
      = ~((~(out_adp_set_value_ac_float_mux_50_nl | (~ operator_5_true_mux_21_nl)))
      | out_adp_set_value_ac_float_lor_11_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_50_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_11_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_11_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_736_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_11_itm_1
      | out_adp_set_value_ac_float_1_mux_90_tmp_3;
  assign operator_5_true_1_mux_21_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_736_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_10_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_50_nl | (~ operator_5_true_1_mux_21_nl)))
      | out_adp_set_value_ac_float_1_lor_11_lpi_1_dfm_1);
  assign write_data_data_10_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_10_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_10_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_10_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign operator_5_true_not_90_nl = ~ NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_43_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_6_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_90_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_43_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_43_nl, 2'b11, out_adp_set_value_ac_float_lor_6_lpi_1_dfm_1));
  assign operator_5_true_1_not_90_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_43_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_6_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_90_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_43_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_43_nl, 2'b11, out_adp_set_value_ac_float_1_lor_6_lpi_1_dfm_1));
  assign write_data_data_5_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_5_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_43_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_43_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_25_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_6_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_6_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_608_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1
      | out_adp_set_value_ac_float_mux_85_tmp_3;
  assign operator_5_true_mux_11_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_608_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_5_nl
      = ~((~(out_adp_set_value_ac_float_mux_25_nl | (~ operator_5_true_mux_11_nl)))
      | out_adp_set_value_ac_float_lor_6_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_25_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_6_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_6_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_706_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1
      | out_adp_set_value_ac_float_1_mux_85_tmp_3;
  assign operator_5_true_1_mux_11_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_706_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_5_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_25_nl | (~ operator_5_true_1_mux_11_nl)))
      | out_adp_set_value_ac_float_1_lor_6_lpi_1_dfm_1);
  assign write_data_data_5_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_5_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_5_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_5_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_15_nl = out_float_round_32_if_m_1_8_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_6_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_15_nl = out_float_round_32_1_if_m_1_8_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_6_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_875_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_5_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_15_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_15_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_27_nl = out_float_round_32_if_m_1_12_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_10_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_27_nl = out_float_round_32_1_if_m_1_12_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_10_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_887_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_9_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_27_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_27_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign operator_5_true_not_98_nl = ~ NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_44_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_10_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_98_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_44_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_44_nl, 2'b11, out_adp_set_value_ac_float_lor_10_lpi_1_dfm_1));
  assign operator_5_true_1_not_98_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_44_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_10_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_98_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_44_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_44_nl, 2'b11, out_adp_set_value_ac_float_1_lor_10_lpi_1_dfm_1));
  assign write_data_data_9_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_9_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_44_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_44_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_45_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_10_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_10_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_632_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1
      | out_adp_set_value_ac_float_mux_89_tmp_3;
  assign operator_5_true_mux_19_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_632_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_9_nl
      = ~((~(out_adp_set_value_ac_float_mux_45_nl | (~ operator_5_true_mux_19_nl)))
      | out_adp_set_value_ac_float_lor_10_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_45_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_10_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_10_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_730_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1
      | out_adp_set_value_ac_float_1_mux_89_tmp_3;
  assign operator_5_true_1_mux_19_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_730_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_9_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_45_nl | (~ operator_5_true_1_mux_19_nl)))
      | out_adp_set_value_ac_float_1_lor_10_lpi_1_dfm_1);
  assign write_data_data_9_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_9_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_9_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_9_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign operator_5_true_not_92_nl = ~ NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_45_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_7_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_92_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_45_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_45_nl, 2'b11, out_adp_set_value_ac_float_lor_7_lpi_1_dfm_1));
  assign operator_5_true_1_not_92_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_45_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_7_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_92_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_45_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_45_nl, 2'b11, out_adp_set_value_ac_float_1_lor_7_lpi_1_dfm_1));
  assign write_data_data_6_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_6_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_45_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_45_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_30_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_7_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_7_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_614_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_7_itm_1
      | out_adp_set_value_ac_float_mux_86_tmp_3;
  assign operator_5_true_mux_13_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_614_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_6_nl
      = ~((~(out_adp_set_value_ac_float_mux_30_nl | (~ operator_5_true_mux_13_nl)))
      | out_adp_set_value_ac_float_lor_7_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_30_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_7_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_7_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_712_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_7_itm_1
      | out_adp_set_value_ac_float_1_mux_86_tmp_3;
  assign operator_5_true_1_mux_13_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_712_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_6_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_30_nl | (~ operator_5_true_1_mux_13_nl)))
      | out_adp_set_value_ac_float_1_lor_7_lpi_1_dfm_1);
  assign write_data_data_6_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_6_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_6_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_6_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_18_nl = out_float_round_32_if_m_1_9_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_7_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_18_nl = out_float_round_32_1_if_m_1_9_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_7_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_878_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_6_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_18_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_18_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_24_nl = out_float_round_32_if_m_1_11_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_9_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_24_nl = out_float_round_32_1_if_m_1_11_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_9_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_884_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_8_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_24_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_24_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign operator_5_true_not_96_nl = ~ NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_46_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_9_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_96_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_46_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_46_nl, 2'b11, out_adp_set_value_ac_float_lor_9_lpi_1_dfm_1));
  assign operator_5_true_1_not_96_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_46_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_9_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_96_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_46_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_46_nl, 2'b11, out_adp_set_value_ac_float_1_lor_9_lpi_1_dfm_1));
  assign write_data_data_8_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_8_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_46_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_46_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_40_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_9_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_9_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_626_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_9_itm_1
      | out_adp_set_value_ac_float_mux_88_tmp_3;
  assign operator_5_true_mux_17_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_626_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_8_nl
      = ~((~(out_adp_set_value_ac_float_mux_40_nl | (~ operator_5_true_mux_17_nl)))
      | out_adp_set_value_ac_float_lor_9_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_40_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_9_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_9_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_724_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_9_itm_1
      | out_adp_set_value_ac_float_1_mux_88_tmp_3;
  assign operator_5_true_1_mux_17_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_724_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_8_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_40_nl | (~ operator_5_true_1_mux_17_nl)))
      | out_adp_set_value_ac_float_1_lor_9_lpi_1_dfm_1);
  assign write_data_data_8_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_8_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_8_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_8_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign operator_5_true_not_94_nl = ~ NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_47_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_exp_tmp_8_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_not_94_nl));
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_47_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_nor_47_nl, 2'b11, out_adp_set_value_ac_float_lor_8_lpi_1_dfm_1));
  assign operator_5_true_1_not_94_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_47_nl = ~(MUX_v_2_2_2((out_adp_set_value_ac_float_1_exp_tmp_8_lpi_1_dfm_4_1_mx0[1:0]),
      2'b11, operator_5_true_1_not_94_nl));
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_47_nl
      = ~(MUX_v_2_2_2(out_adp_set_value_ac_float_1_nor_47_nl, 2'b11, out_adp_set_value_ac_float_1_lor_8_lpi_1_dfm_1));
  assign write_data_data_7_6_4_sva_dfm_1_2_1_mx0w0 = MUX1HOT_v_2_3_2(write_data_data_7_6_4_sva_dfm_1_2_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_47_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_47_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_mux_35_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_acc_sdt_8_sva_1[0]),
      (out_adp_set_value_ac_float_exp_tmp_8_sva_2[0]), NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign or_620_nl = or_dcpl_489 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2) | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1
      | out_adp_set_value_ac_float_mux_87_tmp_3;
  assign operator_5_true_mux_15_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs,
      or_620_nl);
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_7_nl
      = ~((~(out_adp_set_value_ac_float_mux_35_nl | (~ operator_5_true_mux_15_nl)))
      | out_adp_set_value_ac_float_lor_8_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_mux_35_nl = MUX_s_1_2_2((out_adp_set_value_ac_float_1_acc_sdt_8_sva_1[0]),
      (out_adp_set_value_ac_float_1_exp_tmp_8_sva_2[0]), NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign or_718_nl = or_dcpl_587 | NMP_RunFSM_switch_lp_conc_itm_17_2 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1
      | out_adp_set_value_ac_float_1_mux_87_tmp_3;
  assign operator_5_true_1_mux_15_nl = MUX_s_1_2_2(NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0,
      NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs,
      or_718_nl);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_7_nl
      = ~((~(out_adp_set_value_ac_float_1_mux_35_nl | (~ operator_5_true_1_mux_15_nl)))
      | out_adp_set_value_ac_float_1_lor_8_lpi_1_dfm_1);
  assign write_data_data_7_6_4_sva_dfm_1_0_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_7_6_4_sva_dfm_1_0,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_out_adp_set_value_ac_float_nor_7_nl,
      out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_nor_7_nl,
      {while_asn_734 , while_asn_738 , while_asn_740});
  assign out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_21_nl = out_float_round_32_if_m_1_10_sva_1_6
      & (~ out_adp_set_value_ac_float_lor_8_lpi_1_dfm_1);
  assign out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_21_nl = out_float_round_32_1_if_m_1_10_sva_1_6
      & (~ out_adp_set_value_ac_float_1_lor_8_lpi_1_dfm_1);
  assign NMP_RunFSM_switch_lp_mux1h_881_mx0w0 = MUX1HOT_s_1_3_2(write_data_data_7_7_sva_dfm_1,
      out_adp_set_value_ac_float_out_adp_set_value_ac_float_and_21_nl, out_adp_set_value_ac_float_1_out_adp_set_value_ac_float_1_and_21_nl,
      {NMP_RunFSM_switch_lp_or_861_cse_1 , NMP_RunFSM_switch_lp_equal_tmp_4_16 ,
      NMP_RunFSM_switch_lp_equal_tmp_8_16});
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_tmp
      = (NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_1_tmp
      = (NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_2_tmp
      = (NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_3_tmp
      = (NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_4_tmp
      = (NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_5_tmp
      = (NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_6_tmp
      = (NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_7_tmp
      = (NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_8_tmp
      = (NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_9_tmp
      = (NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_10_tmp
      = (NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_11_tmp
      = (NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_12_tmp
      = (NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_13_tmp
      = (NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_14_tmp
      = (NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_15_tmp
      = (NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_out_3[4:1]) < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_1_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_2_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_3_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_4_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_5_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_6_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_7_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_8_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_9_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_10_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_11_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_12_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_13_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_14_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_15_tmp
      = (NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_out_3[4:1])
      < 4'b1101;
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qelse_acc_sdt
      = conv_u2u_39_40(~ (operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp[38:0]))
      + 40'b0000000000000000000000000000000000000001;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qelse_acc_sdt
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qelse_acc_sdt[39:0];
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_mx0_39
      = (ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qelse_acc_sdt[39])
      & (operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp[39]);
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_mx0_38_0
      = MUX_v_39_2_2((operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp[38:0]), (ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qelse_acc_sdt[38:0]),
      operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp[39]);
  assign while_while_while_or_nl = MUX_v_8_2_2(nmp_config_vector_counter_sva_3_1,
      8'b11111111, while_asn_736);
  assign or_922_nl = ((~ mux_cse) & while_asn_736) | NMP_RunFSM_switch_lp_equal_tmp_22
      | NMP_RunFSM_switch_lp_equal_tmp_18_1 | NMP_RunFSM_switch_lp_equal_tmp_20 |
      NMP_RunFSM_switch_lp_equal_tmp_23 | NMP_RunFSM_switch_lp_equal_tmp_17 | NMP_RunFSM_switch_lp_equal_tmp_19
      | NMP_RunFSM_switch_lp_equal_tmp_21 | NMP_RunFSM_switch_lp_equal_tmp_24 | NMP_RunFSM_switch_lp_equal_tmp_25
      | NMP_RunFSM_switch_lp_equal_tmp_10_1 | NMP_RunFSM_switch_lp_equal_tmp_11_1
      | NMP_RunFSM_switch_lp_or_tmp_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign mux_258_nl = MUX_v_8_2_2(while_while_while_or_nl, nmp_config_vector_counter_sva,
      or_922_nl);
  assign nor_266_nl = ~(NMP_RunFSM_switch_lp_and_2_rgt | (mux_cse & while_asn_736));
  assign nmp_config_vector_counter_sva_mx0w0 = MUX_v_8_2_2(8'b00000000, mux_258_nl,
      nor_266_nl);
  assign nmp_config_vector_counter_sva_mx1 = MUX_v_8_2_2(nmp_config_vector_counter_sva,
      nmp_config_vector_counter_sva_mx0w0, while_stage_0_3);
  assign state_3_sva_mx1 = MUX_s_1_2_2(next_state_3_lpi_1_dfm_4, state_3_sva, or_dcpl_481);
  assign state_2_sva_mx1 = MUX_s_1_2_2(next_state_2_lpi_1_dfm_4, state_2_sva, or_dcpl_481);
  assign state_0_sva_mx1 = MUX_s_1_2_2(next_state_0_lpi_1_dfm_4, state_0_sva, or_dcpl_481);
  assign state_1_sva_mx1 = MUX_s_1_2_2(state_1_sva, state_1_sva_dfm_1, while_stage_0_3);
  assign NMP_RunFSM_switch_lp_equal_tmp_13 = state_3_sva_mx1 & state_2_sva_mx1 &
      (~(state_1_sva_mx1 | state_0_sva_mx1));
  assign NMP_RunFSM_switch_lp_equal_tmp_14 = state_1_sva_mx1 & (~(state_3_sva_mx1
      | state_2_sva_mx1 | state_0_sva_mx1));
  assign NMP_RunFSM_switch_lp_equal_tmp_15 = state_3_sva_mx1 & state_1_sva_mx1 &
      state_0_sva_mx1 & (~ state_2_sva_mx1);
  assign NMP_RunFSM_switch_lp_equal_tmp_16 = ~(state_3_sva_mx1 | state_2_sva_mx1
      | state_1_sva_mx1 | state_0_sva_mx1);
  assign NMP_RunFSM_switch_lp_and_2_rgt = (~ nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1)
      & NMP_RunFSM_switch_lp_equal_tmp_12_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nl_operator_8_false_acc_1_nl = 10'b1100000010 + conv_u2s_8_10(~ nmp_config_num_vector_1_sva)
      + conv_u2s_8_10(nmp_config_vector_counter_sva_mx1);
  assign operator_8_false_acc_1_nl = nl_operator_8_false_acc_1_nl[9:0];
  assign operator_8_false_acc_1_itm_9_1 = readslicef_10_1_9(operator_8_false_acc_1_nl);
  assign NMP_UpdateFSM_switch_lp_equal_tmp_7 = state_0_sva_mx1 & (~(state_3_sva_mx1
      | state_2_sva_mx1 | state_1_sva_mx1));
  assign NMP_UpdateFSM_switch_lp_equal_tmp_8 = state_1_sva_mx1 & state_0_sva_mx1
      & (~(state_3_sva_mx1 | state_2_sva_mx1));
  assign NMP_UpdateFSM_switch_lp_equal_tmp_9 = state_2_sva_mx1 & state_1_sva_mx1
      & state_0_sva_mx1 & (~ state_3_sva_mx1);
  assign NMP_UpdateFSM_switch_lp_or_tmp_1_1 = NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_6_cse_1
      | NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_7_cse_1;
  assign NMP_UpdateFSM_switch_lp_nor_tmp_1_1 = ~(NMP_UpdateFSM_switch_lp_equal_tmp_7
      | NMP_UpdateFSM_switch_lp_equal_tmp_8 | NMP_UpdateFSM_switch_lp_equal_tmp_10
      | NMP_UpdateFSM_switch_lp_equal_tmp_11 | NMP_UpdateFSM_switch_lp_equal_tmp_9
      | NMP_UpdateFSM_switch_lp_equal_tmp_12 | NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_6_cse_1
      | NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_7_cse_1 | NMP_UpdateFSM_switch_lp_equal_tmp_13
      | NMP_RunFSM_switch_lp_equal_tmp_15 | NMP_RunFSM_switch_lp_equal_tmp_14 | NMP_RunFSM_switch_lp_equal_tmp_16);
  assign NMP_UpdateFSM_switch_lp_equal_tmp_10 = state_2_sva_mx1 & (~(state_3_sva_mx1
      | state_1_sva_mx1 | state_0_sva_mx1));
  assign NMP_UpdateFSM_switch_lp_equal_tmp_11 = state_2_sva_mx1 & state_1_sva_mx1
      & (~(state_3_sva_mx1 | state_0_sva_mx1));
  assign NMP_UpdateFSM_switch_lp_equal_tmp_12 = state_3_sva_mx1 & (~(state_2_sva_mx1
      | state_1_sva_mx1 | state_0_sva_mx1));
  assign NMP_UpdateFSM_switch_lp_equal_tmp_13 = state_3_sva_mx1 & state_1_sva_mx1
      & (~(state_2_sva_mx1 | state_0_sva_mx1));
  assign nl_out_adp_set_value_ac_float_acc_sdt_1_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_1_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_1_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_1_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_2_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_1_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_2_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_2_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_2_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_3_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_2_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_3_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_3_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_3_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_4_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_3_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_4_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_4_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_4_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_5_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_4_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_5_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_5_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_5_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_6_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_5_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_6_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_6_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_6_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_7_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_6_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_7_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_7_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_7_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_8_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_7_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_8_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_8_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_8_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_9_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_8_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_9_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_9_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_9_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_10_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_9_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_10_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_10_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_10_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_11_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_10_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_11_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_11_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_11_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_12_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_11_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_12_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_12_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_12_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_13_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_12_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_13_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_13_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_13_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_14_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_13_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_14_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_14_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_14_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_15_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_14_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_15_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_15_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_15_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_acc_sdt_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_15_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_acc_sdt_sva_1 = nl_out_adp_set_value_ac_float_acc_sdt_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_exp_tmp_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_1_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_1_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_1_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_1_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_2_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_1_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_2_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_2_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_2_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_3_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_2_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_3_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_3_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_3_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_4_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_3_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_4_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_4_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_4_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_5_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_4_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_5_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_5_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_5_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_6_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_5_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_6_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_6_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_6_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_7_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_6_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_7_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_7_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_7_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_8_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_7_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_8_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_8_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_8_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_9_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_8_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_9_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_9_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_9_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_10_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_9_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_10_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_10_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_10_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_11_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_10_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_11_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_11_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_11_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_12_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_11_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_12_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_12_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_12_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_13_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_12_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_13_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_13_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_13_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_14_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_13_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_14_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_14_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_14_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_15_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_14_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_15_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_15_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_15_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_out_adp_set_value_ac_float_1_acc_sdt_sva_1 = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_15_itm_1
      + conv_s2u_4_5({1'b1 , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd)
      , (~ reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1)}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_acc_sdt_sva_1 = nl_out_adp_set_value_ac_float_1_acc_sdt_sva_1[4:0];
  assign NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0
      = ~((out_adp_set_value_ac_float_1_exp_tmp_lpi_1_dfm_4_1_mx0[3:2]==2'b01));
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_mx0w0
      = $signed(({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_itm}))
      * $signed(conv_u2s_10_11(ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_itm));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_mx0w0
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_mx0w0[18:0];
  assign NMP_RunFSM_switch_lp_and_24_nl = (~ NMP_ComputeSoftmaxMax_for_if_slc_NMP_ComputeSoftmaxMax_for_16_acc_1_27_svs_1)
      & NMP_RunFSM_switch_lp_equal_tmp_5_4;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux1h_3_nl = MUX1HOT_s_1_3_2(max_value_26_0_sva_26,
      max_value_26_0_sva_dfm_14_26_mx0, (reg_NMP_RunFSM_switch_lp_asn_104_itm_3_cse[26]),
      {(~ NMP_RunFSM_switch_lp_equal_tmp_5_4) , NMP_RunFSM_switch_lp_and_24_nl ,
      NMP_RunFSM_switch_lp_and_25_ssc_1});
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_54_itm = NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux1h_3_nl
      & (~ NMP_RunFSM_switch_lp_equal_tmp_5);
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux_2_nl
      = MUX_v_26_2_2(max_value_26_0_sva_dfm_14_25_0_mx0, (reg_NMP_RunFSM_switch_lp_asn_104_itm_3_cse[25:0]),
      NMP_RunFSM_switch_lp_and_25_ssc_1);
  assign NMP_RunFSM_switch_lp_not_80_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_5;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_52_itm = MUX_v_26_2_2(26'b00000000000000000000000000,
      NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_mux_2_nl, NMP_RunFSM_switch_lp_not_80_nl);
  assign or_924_itm = (~(NMP_RunFSM_switch_lp_equal_tmp_5 | NMP_RunFSM_switch_lp_equal_tmp_5_4))
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign NMP_RunFSM_switch_lp_and_25_ssc_1 = NMP_ComputeSoftmaxMax_for_if_slc_NMP_ComputeSoftmaxMax_for_16_acc_1_27_svs_1
      & NMP_RunFSM_switch_lp_equal_tmp_5_4;
  assign nmp_config_adpbias_1_sva_mx1_2 = MUX_s_1_2_2(reg_nmp_config_adpbias_1_ftd,
      nmp_config_adpbias_1_sva_dfm_3_1_2, while_stage_0_3);
  assign nmp_config_adpbias_1_sva_mx1_1_0 = MUX_v_2_2_2(reg_nmp_config_adpbias_1_ftd_1,
      nmp_config_adpbias_1_sva_dfm_3_1_1_0, while_stage_0_3);
  assign nl_sum_exp_39_4_sva_1 = conv_u2u_34_36(NMP_ComputeSoftmaxSum_for_acc_7_itm_1)
      + conv_u2u_34_36(NMP_ComputeSoftmaxSum_for_acc_8_itm_1) + conv_u2u_34_36(NMP_ComputeSoftmaxSum_for_acc_9_itm_1)
      + conv_u2u_34_36(NMP_ComputeSoftmaxSum_for_acc_11_itm_1) + conv_u2u_33_36(NMP_ComputeSoftmaxSum_for_acc_12_itm_1)
      + conv_u2u_33_36(NMP_ComputeSoftmaxSum_for_acc_13_itm_1);
  assign sum_exp_39_4_sva_1 = nl_sum_exp_39_4_sva_1[35:0];
  assign max_value_26_0_sva_dfm_9_1_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_8_26_mx0,
      (NMP_ComputeSoftmaxExp_for_asn_24_itm_1[26]), NMP_ComputeSoftmaxMax_for_if_less_6_itm);
  assign NMP_ComputeSoftmaxMax_for_if_less_5_tmp = $signed(({max_value_26_0_sva_dfm_9_1_26_mx0
      , max_value_26_0_sva_dfm_9_1_25_0_mx0})) < $signed(NMP_ComputeSoftmaxExp_for_asn_25_itm_1);
  assign max_value_26_0_sva_dfm_9_1_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_8_25_0_mx0,
      (NMP_ComputeSoftmaxExp_for_asn_24_itm_1[25:0]), NMP_ComputeSoftmaxMax_for_if_less_6_itm);
  assign NMP_RunFSM_switch_lp_not_81_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_31_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_16_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_81_nl);
  assign exp_values_15_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_31_nl,
      exp_values_15_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_82_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_30_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_15_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_82_nl);
  assign exp_values_14_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_30_nl,
      exp_values_14_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_83_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_29_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_14_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_83_nl);
  assign exp_values_13_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_29_nl,
      exp_values_13_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_84_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_28_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_13_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_84_nl);
  assign exp_values_12_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_28_nl,
      exp_values_12_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_85_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_27_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_12_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_85_nl);
  assign exp_values_11_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_27_nl,
      exp_values_11_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_86_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_26_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_11_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_86_nl);
  assign exp_values_10_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_26_nl,
      exp_values_10_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_87_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_25_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_10_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_87_nl);
  assign exp_values_9_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_25_nl,
      exp_values_9_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_88_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_24_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_9_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_88_nl);
  assign exp_values_8_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_24_nl,
      exp_values_8_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_89_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_23_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_8_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_89_nl);
  assign exp_values_7_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_23_nl,
      exp_values_7_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_90_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_22_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_7_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_90_nl);
  assign exp_values_6_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_22_nl,
      exp_values_6_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_91_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_21_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_6_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_91_nl);
  assign exp_values_5_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_21_nl,
      exp_values_5_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_92_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_20_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_5_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_92_nl);
  assign exp_values_4_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_20_nl,
      exp_values_4_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_93_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_19_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_4_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_93_nl);
  assign exp_values_3_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_19_nl,
      exp_values_3_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_94_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_18_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_3_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_94_nl);
  assign exp_values_2_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_18_nl,
      exp_values_2_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_95_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_17_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_2_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_95_nl);
  assign exp_values_1_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_17_nl,
      exp_values_1_sva, or_dcpl_742);
  assign NMP_RunFSM_switch_lp_not_57_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_8;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_55_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      NMP_ComputeSoftmaxExp_for_1_operator_32_12_false_AC_TRN_AC_WRAP_lshift_itm,
      NMP_RunFSM_switch_lp_not_57_nl);
  assign exp_values_0_sva_mx1 = MUX_v_32_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_55_nl,
      exp_values_0_sva, or_dcpl_742);
  assign nmp_config_mode_sva_mx1 = MUX_v_3_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[3:1]),
      nmp_config_mode_sva, or_dcpl_480);
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_2
      = (operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp!=40'b0000000000000000000000000000000000000000);
  assign max_value_26_0_sva_dfm_2_1_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_1_26_1,
      (input_fixed_2_26_0_sva[26]), NMP_ComputeSoftmaxMax_for_if_less_13_itm);
  assign NMP_ComputeSoftmaxMax_for_if_less_12_tmp = $signed(({max_value_26_0_sva_dfm_2_1_26_mx0
      , max_value_26_0_sva_dfm_2_1_25_0_mx0})) < $signed(input_fixed_mux_9_cse);
  assign max_value_26_0_sva_dfm_2_1_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_1_25_0_mx0,
      (input_fixed_2_26_0_sva[25:0]), NMP_ComputeSoftmaxMax_for_if_less_13_itm);
  assign NMP_RunFSM_switch_lp_equal_tmp_17 = state_2_sva & state_1_sva & (~(state_3_sva
      | state_0_sva));
  assign NMP_RunFSM_switch_lp_not_25_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_4;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_35_nl = MUX_v_36_2_2(36'b000000000000000000000000000000000000,
      sum_sq_1_39_4_sva_2_1, NMP_RunFSM_switch_lp_not_25_nl);
  assign or_927_nl = (~(NMP_RunFSM_switch_lp_equal_tmp_4 | NMP_RunFSM_switch_lp_equal_tmp_2_3))
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ while_stage_0_6);
  assign sum_sq_1_39_4_sva_mx1 = MUX_v_36_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_35_nl,
      sum_sq_1_39_4_sva, or_927_nl);
  assign NMP_RunFSM_switch_lp_equal_tmp_18_1 = state_1_sva & state_0_sva & (~(state_3_sva
      | state_2_sva));
  assign NMP_RunFSM_switch_lp_equal_tmp_19 = state_2_sva & state_1_sva & state_0_sva
      & (~ state_3_sva);
  assign NMP_RunFSM_switch_lp_equal_tmp_20 = state_2_sva & (~(state_3_sva | state_1_sva
      | state_0_sva));
  assign NMP_RunFSM_switch_lp_equal_tmp_21 = state_3_sva & (~(state_2_sva | state_1_sva
      | state_0_sva));
  assign NMP_RunFSM_switch_lp_equal_tmp_22 = state_0_sva & (~(state_3_sva | state_2_sva
      | state_1_sva));
  assign NMP_RunFSM_switch_lp_equal_tmp_23 = state_2_sva & state_0_sva & (~(state_3_sva
      | state_1_sva));
  assign NMP_RunFSM_switch_lp_equal_tmp_24 = state_3_sva & state_0_sva & (~(state_2_sva
      | state_1_sva));
  assign NMP_RunFSM_switch_lp_equal_tmp_25 = state_3_sva & state_1_sva & (~(state_2_sva
      | state_0_sva));
  assign NMP_RunFSM_switch_lp_or_tmp_1 = (state_3_sva & state_2_sva & state_0_sva
      & (~ state_1_sva)) | (state_3_sva & state_2_sva & state_1_sva & (~ state_0_sva))
      | (state_3_sva & state_2_sva & state_1_sva & state_0_sva);
  assign nl_out_adp_set_value_ac_float_exp_tmp_1_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_1_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_1_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_1_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_1_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_1_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_1_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_1_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_1_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_1_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_1_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_1_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_2_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_2_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_2_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_2_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_2_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_2_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_2_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_2_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_2_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_2_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_2_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_2_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_3_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_3_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_3_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_3_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_3_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_3_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_3_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_3_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_3_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_3_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_3_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_3_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_4_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_4_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_4_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_4_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_4_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_4_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_4_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_4_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_4_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_4_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_4_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_4_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_5_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_5_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_5_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_5_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_5_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_5_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_5_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_5_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_5_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_5_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_5_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_5_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_6_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_6_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_6_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_6_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_6_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_6_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_6_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_6_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_6_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_6_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_6_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_6_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_7_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_7_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_7_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_7_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_7_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_7_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_7_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_7_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_7_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_7_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_7_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_7_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_8_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_8_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_8_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_8_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_8_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_8_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_8_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_8_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_8_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_8_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_8_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_8_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_9_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_9_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_9_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_9_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_9_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_9_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_9_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_9_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_9_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_9_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_9_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_9_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_10_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_10_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_10_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_10_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_10_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_10_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_10_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_10_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_10_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_10_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_10_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_10_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_11_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_11_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_11_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_11_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_11_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_11_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_11_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_11_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_11_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_11_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_11_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_11_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_12_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_12_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_12_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_12_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_12_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_12_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_12_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_12_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_12_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_12_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_12_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_12_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_13_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_13_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_13_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_13_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_13_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_13_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_13_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_13_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_13_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_13_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_13_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_13_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_14_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_14_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_14_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_14_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_14_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_14_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_14_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_14_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_14_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_14_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_14_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_14_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_15_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_15_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_15_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_15_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_15_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_15_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_15_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_15_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_15_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_15_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_15_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_15_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign nl_out_adp_set_value_ac_float_exp_tmp_sva_2 = ({out_adp_set_value_ac_float_ac_int_cctor_4_1_sva_1
      , (out_adp_set_value_ac_float_acc_sdt_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_exp_tmp_sva_2 = nl_out_adp_set_value_ac_float_exp_tmp_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_acc_sdt_sva_1[4:1]);
  assign out_adp_set_value_ac_float_ac_int_cctor_4_1_sva_1 = nl_out_adp_set_value_ac_float_ac_int_cctor_4_1_sva_1[3:0];
  assign out_adp_set_value_ac_float_exp_tmp_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_ac_int_cctor_4_1_sva_1,
      (out_adp_set_value_ac_float_exp_tmp_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_lor_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_16_itm_1;
  assign out_adp_set_value_ac_float_lor_15_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_15_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1;
  assign out_adp_set_value_ac_float_lor_14_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_14_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_14_itm_1;
  assign out_adp_set_value_ac_float_lor_13_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_13_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_13_itm_1;
  assign out_adp_set_value_ac_float_lor_12_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_12_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1;
  assign out_adp_set_value_ac_float_lor_11_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_11_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1;
  assign out_adp_set_value_ac_float_lor_10_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_10_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1;
  assign out_adp_set_value_ac_float_lor_9_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_9_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_9_itm_1;
  assign out_adp_set_value_ac_float_lor_8_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_8_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1;
  assign out_adp_set_value_ac_float_lor_7_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_7_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_7_itm_1;
  assign out_adp_set_value_ac_float_lor_6_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_6_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1;
  assign out_adp_set_value_ac_float_lor_5_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_5_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1;
  assign out_adp_set_value_ac_float_lor_4_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_4_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_4_itm_1;
  assign out_adp_set_value_ac_float_lor_3_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_3_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_3_itm_1;
  assign out_adp_set_value_ac_float_lor_2_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_2_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_2_itm_1;
  assign out_adp_set_value_ac_float_lor_1_lpi_1_dfm_1 = (out_adp_set_value_ac_float_exp_tmp_1_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_itm_1;
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_1_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_1_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_1_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_1_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_1_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_1_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_1_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_1_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_1_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_1_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_1_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_1_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_2_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_2_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_2_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_2_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_2_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_2_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_2_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_2_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_2_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_2_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_2_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_2_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_3_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_3_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_3_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_3_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_3_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_3_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_3_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_3_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_3_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_3_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_3_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_3_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_4_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_4_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_4_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_4_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_4_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_4_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_4_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_4_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_4_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_4_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_4_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_4_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_5_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_5_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_5_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_5_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_5_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_5_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_5_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_5_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_5_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_5_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_5_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_5_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_6_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_6_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_6_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_6_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_6_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_6_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_6_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_6_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_6_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_6_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_6_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_6_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_7_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_7_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_7_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_7_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_7_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_7_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_7_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_7_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_7_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_7_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_7_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_7_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_8_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_8_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_8_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_8_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_8_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_8_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_8_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_8_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_8_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_8_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_8_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_8_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_9_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_9_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_9_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_9_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_9_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_9_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_9_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_9_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_9_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_9_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_9_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_9_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_10_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_10_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_10_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_10_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_10_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_10_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_10_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_10_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_10_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_10_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_10_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_10_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_11_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_11_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_11_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_11_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_11_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_11_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_11_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_11_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_11_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_11_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_11_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_11_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_12_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_12_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_12_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_12_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_12_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_12_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_12_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_12_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_12_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_12_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_12_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_12_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_13_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_13_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_13_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_13_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_13_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_13_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_13_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_13_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_13_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_13_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_13_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_13_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_14_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_14_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_14_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_14_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_14_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_14_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_14_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_14_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_14_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_14_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_14_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_14_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_15_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_15_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_15_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_15_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_15_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_15_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_15_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_15_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_15_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_15_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_15_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_15_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign nl_out_adp_set_value_ac_float_1_exp_tmp_sva_2 = ({out_adp_set_value_ac_float_1_ac_int_cctor_4_1_sva_1
      , (out_adp_set_value_ac_float_1_acc_sdt_sva_1[0])}) + 5'b00001;
  assign out_adp_set_value_ac_float_1_exp_tmp_sva_2 = nl_out_adp_set_value_ac_float_1_exp_tmp_sva_2[4:0];
  assign nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_sva_1 = 4'b0101 + (out_adp_set_value_ac_float_1_acc_sdt_sva_1[4:1]);
  assign out_adp_set_value_ac_float_1_ac_int_cctor_4_1_sva_1 = nl_out_adp_set_value_ac_float_1_ac_int_cctor_4_1_sva_1[3:0];
  assign out_adp_set_value_ac_float_1_exp_tmp_lpi_1_dfm_4_1_mx0 = MUX_v_4_2_2(out_adp_set_value_ac_float_1_ac_int_cctor_4_1_sva_1,
      (out_adp_set_value_ac_float_1_exp_tmp_sva_2[4:1]), NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_lor_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_16_itm_1;
  assign out_adp_set_value_ac_float_1_lor_15_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_15_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_15_itm_1;
  assign out_adp_set_value_ac_float_1_lor_14_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_14_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1;
  assign out_adp_set_value_ac_float_1_lor_13_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_13_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_13_itm_1;
  assign out_adp_set_value_ac_float_1_lor_12_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_12_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_12_itm_1;
  assign out_adp_set_value_ac_float_1_lor_11_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_11_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_11_itm_1;
  assign out_adp_set_value_ac_float_1_lor_10_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_10_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1;
  assign out_adp_set_value_ac_float_1_lor_9_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_9_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_9_itm_1;
  assign out_adp_set_value_ac_float_1_lor_8_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_8_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1;
  assign out_adp_set_value_ac_float_1_lor_7_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_7_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_7_itm_1;
  assign out_adp_set_value_ac_float_1_lor_6_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_6_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1;
  assign out_adp_set_value_ac_float_1_lor_5_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_5_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_5_itm_1;
  assign out_adp_set_value_ac_float_1_lor_4_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_4_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1;
  assign out_adp_set_value_ac_float_1_lor_3_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_3_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1;
  assign out_adp_set_value_ac_float_1_lor_2_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_2_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1;
  assign out_adp_set_value_ac_float_1_lor_1_lpi_1_dfm_1 = (out_adp_set_value_ac_float_1_exp_tmp_1_lpi_1_dfm_4_1_mx0[3])
      | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1;
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_qif_ac_fixed_cctor_20_0_sva_1
      = ({(~ ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_psp_sva)
      , (~ ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1_9_0)})
      + 21'b000000000000000000001;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_qif_ac_fixed_cctor_20_0_sva_1
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_1_if_qif_ac_fixed_cctor_20_0_sva_1[20:0];
  assign NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_25_nl = (~ NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2)
      & large_rsp_PopNB_mioi_return_rsc_z_mxwt;
  assign NMP_RunFSM_switch_lp_mux1h_74_nl = MUX1HOT_s_1_4_2(mux_cse, state_0_sva,
      NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_25_nl, (~ NMP_UpdateFSM_case_11_time_end_lpi_1_dfm_1),
      {NMP_RunFSM_switch_lp_equal_tmp_1 , NMP_RunFSM_switch_lp_or_73_tmp , NMP_RunFSM_switch_lp_equal_tmp_11_1
      , NMP_RunFSM_switch_lp_equal_tmp_12_1});
  assign next_state_0_lpi_1_dfm_4 = (NMP_RunFSM_switch_lp_mux1h_74_nl & (~(NMP_UpdateFSM_switch_lp_equal_tmp_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_1_1 | NMP_UpdateFSM_switch_lp_equal_tmp_4_1
      | NMP_UpdateFSM_switch_lp_or_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1))) |
      NMP_UpdateFSM_switch_lp_equal_tmp_2_1 | NMP_UpdateFSM_switch_lp_equal_tmp_3_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_5_1 | NMP_UpdateFSM_switch_lp_equal_tmp_6_1;
  assign NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_24_nl = NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2
      & large_rsp_PopNB_mioi_return_rsc_z_mxwt;
  assign NMP_RunFSM_switch_lp_mux1h_72_nl = MUX1HOT_s_1_3_2(state_2_sva, NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_24_nl,
      NMP_UpdateFSM_case_11_time_end_lpi_1_dfm_1, {NMP_RunFSM_switch_lp_or_73_tmp
      , NMP_RunFSM_switch_lp_equal_tmp_11_1 , NMP_RunFSM_switch_lp_equal_tmp_12_1});
  assign next_state_2_lpi_1_dfm_4 = (NMP_RunFSM_switch_lp_mux1h_72_nl & (~ NMP_RunFSM_switch_lp_equal_tmp_1)
      & (~(NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_equal_tmp_4_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_5_1 | NMP_UpdateFSM_switch_lp_or_tmp_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_6_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1)))
      | NMP_UpdateFSM_switch_lp_equal_tmp_1_1 | NMP_UpdateFSM_switch_lp_equal_tmp_2_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_3_1;
  assign NMP_RunFSM_switch_lp_mux_51_nl = MUX_s_1_2_2(next_state_3_lpi_1_dfm_3, NMP_UpdateFSM_case_11_time_end_lpi_1_dfm_1,
      NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign next_state_3_lpi_1_dfm_4 = (NMP_RunFSM_switch_lp_mux_51_nl & (~ NMP_RunFSM_switch_lp_equal_tmp_11_1)
      & (~ NMP_RunFSM_switch_lp_equal_tmp_1) & (~(NMP_UpdateFSM_switch_lp_equal_tmp_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_1_1 | NMP_UpdateFSM_switch_lp_equal_tmp_2_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_3_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1)))
      | NMP_UpdateFSM_switch_lp_equal_tmp_4_1 | NMP_UpdateFSM_switch_lp_equal_tmp_5_1
      | NMP_UpdateFSM_switch_lp_or_tmp_1 | NMP_UpdateFSM_switch_lp_equal_tmp_6_1;
  assign in_adp_is_zero_land_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[126:120]!=7'b0000000));
  assign in_adp_is_zero_land_15_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[118:112]!=7'b0000000));
  assign in_adp_is_zero_land_14_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[110:104]!=7'b0000000));
  assign in_adp_is_zero_land_13_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[102:96]!=7'b0000000));
  assign in_adp_is_zero_land_12_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[94:88]!=7'b0000000));
  assign in_adp_is_zero_land_11_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[86:80]!=7'b0000000));
  assign in_adp_is_zero_land_10_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[78:72]!=7'b0000000));
  assign in_adp_is_zero_land_9_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[70:64]!=7'b0000000));
  assign in_adp_is_zero_land_8_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[62:56]!=7'b0000000));
  assign in_adp_is_zero_land_7_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[54:48]!=7'b0000000));
  assign in_adp_is_zero_land_6_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[46:40]!=7'b0000000));
  assign in_adp_is_zero_land_5_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[38:32]!=7'b0000000));
  assign in_adp_is_zero_land_4_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[30:24]!=7'b0000000));
  assign in_adp_is_zero_land_3_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[22:16]!=7'b0000000));
  assign in_adp_is_zero_land_2_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[14:8]!=7'b0000000));
  assign in_adp_is_zero_land_1_lpi_1_dfm_1 = ~((large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[6:0]!=7'b0000000));
  assign NMP_UpdateFSM_case_11_time_end_lpi_1_dfm_1 = ~(operator_16_false_acc_2_itm_17
      | nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1);
  assign nl_operator_16_false_acc_2_nl_1 = 18'b110000000000000010 + conv_u2s_16_18(~
      nmp_config_num_timestep_1_sva) + conv_u2s_16_18(nmp_config_timestep_counter_sva);
  assign operator_16_false_acc_2_nl_1 = nl_operator_16_false_acc_2_nl_1[17:0];
  assign operator_16_false_acc_2_itm_17 = readslicef_18_1_17(operator_16_false_acc_2_nl_1);
  assign NMP_RunFSM_switch_lp_or_73_tmp = NMP_RunFSM_switch_lp_equal_tmp_22 | NMP_RunFSM_switch_lp_equal_tmp_18_1
      | NMP_RunFSM_switch_lp_equal_tmp_20 | NMP_RunFSM_switch_lp_equal_tmp_23 | NMP_RunFSM_switch_lp_equal_tmp_17
      | NMP_RunFSM_switch_lp_equal_tmp_19 | NMP_RunFSM_switch_lp_equal_tmp_21 | NMP_RunFSM_switch_lp_equal_tmp_24
      | NMP_RunFSM_switch_lp_equal_tmp_25 | NMP_RunFSM_switch_lp_equal_tmp_10_1 |
      NMP_RunFSM_switch_lp_or_tmp_1;
  assign NMP_RunFSM_switch_lp_or_861_cse_1 = NMP_RunFSM_switch_lp_equal_tmp_17_1
      | NMP_RunFSM_switch_lp_equal_tmp_1_16 | NMP_RunFSM_switch_lp_equal_tmp_2_16
      | NMP_RunFSM_switch_lp_equal_tmp_3_16 | NMP_RunFSM_switch_lp_equal_tmp_5_16
      | NMP_RunFSM_switch_lp_equal_tmp_6_16 | NMP_RunFSM_switch_lp_equal_tmp_7_16
      | NMP_RunFSM_switch_lp_equal_tmp_9_16 | NMP_RunFSM_switch_lp_equal_tmp_10_17
      | NMP_RunFSM_switch_lp_equal_tmp_11_17 | NMP_RunFSM_switch_lp_equal_tmp_12_17
      | NMP_RunFSM_switch_lp_or_tmp_16;
  assign nl_NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_16_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_16_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_15_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_15_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_14_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_14_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_13_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_13_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_12_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_12_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_11_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_11_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_10_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_10_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp =
      conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_9_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_9_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp =
      conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_8_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_8_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp =
      conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_7_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_7_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp =
      conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_6_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_6_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp =
      conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_5_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_5_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp =
      conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_4_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_4_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp =
      conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_3_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_3_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp =
      conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_2_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_2_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp =
      conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_for_1_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_for_1_operator_32_12_true_AC_TRN_AC_WRAP_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp = nl_NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_16_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_16_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_15_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_15_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_14_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_14_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_13_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_13_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_12_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_12_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_11_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_11_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_10_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_10_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_9_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_9_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_8_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_8_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_7_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_7_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_6_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_6_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_5_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_5_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_4_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_4_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_3_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_3_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_2_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_2_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp
      = conv_s2u_6_7(NMP_ConvertOutputToAdpfloat_1_for_1_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[31:26])
      + conv_u2u_1_7(NMP_ConvertOutputToAdpfloat_1_for_1_operator_32_12_true_AC_TRN_AC_WRAP_1_lshift_itm[25]);
  assign NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp
      = nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp[6:0];
  assign out_float_round_32_rnd_ovfl_1_sva_1 = (NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_2_sva_1 = (NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_3_sva_1 = (NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_4_sva_1 = (NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_5_sva_1 = (NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_6_sva_1 = (NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_7_sva_1 = (NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_8_sva_1 = (NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_9_sva_1 = (NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_10_sva_1 = (NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_11_sva_1 = (NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_12_sva_1 = (NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_13_sva_1 = (NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_14_sva_1 = (NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_15_sva_1 = (NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_rnd_ovfl_sva_1 = (NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp[6:5]==2'b01);
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_sva_1 = (NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_15_sva_1 = (NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_15_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_14_sva_1 = (NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_14_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_13_sva_1 = (NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_13_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_12_sva_1 = (NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_12_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_11_sva_1 = (NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_11_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_10_sva_1 = (NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_10_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_9_sva_1 = (NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_9_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_8_sva_1 = (NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_8_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_7_sva_1 = (NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_7_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_6_sva_1 = (NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_6_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_5_sva_1 = (NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_5_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_4_sva_1 = (NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_4_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_3_sva_1 = (NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_3_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_2_sva_1 = (NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_2_sva_1;
  assign NMP_ConvertOutputToAdpfloat_for_out_float_m_4_1_sva_1 = (NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp[4])
      | out_float_round_32_rnd_ovfl_1_sva_1;
  assign out_float_round_32_1_rnd_ovfl_1_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_2_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_3_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_4_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_5_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_6_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_7_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_8_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_9_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_10_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_11_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_12_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_13_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_14_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_15_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign out_float_round_32_1_rnd_ovfl_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp[6:5]==2'b01);
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_15_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_15_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_14_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_14_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_13_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_13_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_12_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_12_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_11_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_11_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_10_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_10_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_9_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_9_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_8_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_8_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_7_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_7_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_6_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_6_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_5_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_5_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_4_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_4_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_3_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_3_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_2_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_2_sva_1;
  assign NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_1_sva_1 = (NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp[4])
      | out_float_round_32_1_rnd_ovfl_1_sva_1;
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = $signed(({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_itm}))
      * $signed(conv_u2s_10_11(ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_itm));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:0];
  assign nl_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_nl
      = 13'b1011010100001 * ({ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_12_9
      , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_8_0
      , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_7
      , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_6_0});
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_nl
      = nl_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_nl[35:0];
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_itm_35_11_1
      = readslicef_36_25_11(ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_nl);
  assign max_value_26_0_sva_dfm_14_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_13_1_26,
      (NMP_ComputeSoftmaxMax_for_asn_13_itm_3[26]), NMP_ComputeSoftmaxMax_for_if_less_1_itm);
  assign max_value_26_0_sva_dfm_14_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_13_1_25_0,
      (NMP_ComputeSoftmaxMax_for_asn_13_itm_3[25:0]), NMP_ComputeSoftmaxMax_for_if_less_1_itm);
  assign NMP_ComputeSoftmaxMax_for_if_slc_NMP_ComputeSoftmaxMax_for_16_acc_1_27_svs_1
      = $signed(({max_value_26_0_sva_dfm_14_26_mx0 , max_value_26_0_sva_dfm_14_25_0_mx0}))
      < $signed(reg_NMP_RunFSM_switch_lp_asn_104_itm_3_cse);
  assign nmp_config_ConfigRead_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
      & nmp_config_ConfigRead_nor_2_tmp);
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_1_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[3:0]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_1_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_1_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_1_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[6:4])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_1_sva_1 = nl_in_adp_to_ac_float_acc_sdt_1_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_2_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[11:8]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_2_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_2_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_2_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[14:12])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_2_sva_1 = nl_in_adp_to_ac_float_acc_sdt_2_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_3_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[19:16]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_3_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_3_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_3_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[22:20])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_3_sva_1 = nl_in_adp_to_ac_float_acc_sdt_3_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_4_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[27:24]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_4_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_4_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_4_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[30:28])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_4_sva_1 = nl_in_adp_to_ac_float_acc_sdt_4_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_5_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[35:32]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_5_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_5_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_5_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[38:36])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_5_sva_1 = nl_in_adp_to_ac_float_acc_sdt_5_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_6_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[43:40]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_6_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_6_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_6_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[46:44])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_6_sva_1 = nl_in_adp_to_ac_float_acc_sdt_6_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_7_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[51:48]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_7_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_7_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_7_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[54:52])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_7_sva_1 = nl_in_adp_to_ac_float_acc_sdt_7_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_8_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[59:56]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_8_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_8_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_8_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[62:60])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_8_sva_1 = nl_in_adp_to_ac_float_acc_sdt_8_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_9_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[67:64]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_9_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_9_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_9_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[70:68])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_9_sva_1 = nl_in_adp_to_ac_float_acc_sdt_9_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_10_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[75:72]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_10_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_10_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_10_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[78:76])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_10_sva_1 = nl_in_adp_to_ac_float_acc_sdt_10_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_11_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[83:80]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_11_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_11_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_11_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[86:84])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_11_sva_1 = nl_in_adp_to_ac_float_acc_sdt_11_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_12_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[91:88]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_12_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_12_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_12_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[94:92])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_12_sva_1 = nl_in_adp_to_ac_float_acc_sdt_12_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_13_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[99:96]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_13_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_13_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_13_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[102:100])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_13_sva_1 = nl_in_adp_to_ac_float_acc_sdt_13_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_14_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[107:104]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_14_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_14_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_14_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[110:108])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_14_sva_1 = nl_in_adp_to_ac_float_acc_sdt_14_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_15_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[115:112]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_15_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_15_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_15_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[118:116])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_15_sva_1 = nl_in_adp_to_ac_float_acc_sdt_15_sva_1[3:0];
  assign nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_sva_1 = conv_u2s_4_5(~ (large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[123:120]))
      + 5'b00001;
  assign in_adp_to_ac_float_if_1_ac_int_cctor_4_0_sva_1 = nl_in_adp_to_ac_float_if_1_ac_int_cctor_4_0_sva_1[4:0];
  assign nl_in_adp_to_ac_float_acc_sdt_sva_1 = conv_u2u_3_4(large_rsp_PopNB_mioi_data_read_vector_data_data_rsc_z_mxwt[126:124])
      + conv_u2u_3_4({reg_nmp_config_adpbias_1_ftd , reg_nmp_config_adpbias_1_ftd_1});
  assign in_adp_to_ac_float_acc_sdt_sva_1 = nl_in_adp_to_ac_float_acc_sdt_sva_1[3:0];
  assign NMP_RunFSM_switch_lp_and_8_cse_1 = large_rsp_PopNB_mioi_return_rsc_z_mxwt
      & NMP_RunFSM_switch_lp_equal_tmp_11_1;
  assign next_state_1_lpi_1_dfm_4 = ((next_state_1_lpi_1_dfm_3 | NMP_RunFSM_switch_lp_equal_tmp_14)
      & (~(NMP_RunFSM_switch_lp_equal_tmp_16 | NMP_RunFSM_switch_lp_equal_tmp_15))
      & (~(NMP_UpdateFSM_switch_lp_equal_tmp_8 | NMP_UpdateFSM_switch_lp_equal_tmp_10
      | NMP_UpdateFSM_switch_lp_equal_tmp_9 | NMP_UpdateFSM_switch_lp_equal_tmp_12
      | NMP_UpdateFSM_switch_lp_nor_tmp_1_1))) | NMP_UpdateFSM_switch_lp_equal_tmp_7
      | NMP_UpdateFSM_switch_lp_equal_tmp_11 | NMP_UpdateFSM_switch_lp_or_tmp_1_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_13;
  assign NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_6_cse_1 = state_3_sva_mx1
      & state_0_sva_mx1 & (~(state_2_sva_mx1 | state_1_sva_mx1));
  assign NMP_UpdateFSM_switch_lp_NMP_UpdateFSM_switch_lp_and_7_cse_1 = state_2_sva_mx1
      & state_0_sva_mx1 & (~(state_3_sva_mx1 | state_1_sva_mx1));
  assign max_value_26_0_sva_dfm_12_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_11_26_mx0,
      (NMP_ComputeSoftmaxExp_for_asn_27_itm_2[26]), NMP_ComputeSoftmaxMax_for_if_less_3_itm);
  assign max_value_26_0_sva_dfm_12_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_11_25_0_mx0,
      (NMP_ComputeSoftmaxExp_for_asn_27_itm_2[25:0]), NMP_ComputeSoftmaxMax_for_if_less_3_itm);
  assign max_value_26_0_sva_dfm_11_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_10_26_mx0,
      (NMP_ComputeSoftmaxExp_for_asn_26_itm_2[26]), NMP_ComputeSoftmaxMax_for_if_less_4_itm);
  assign max_value_26_0_sva_dfm_11_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_10_25_0_mx0,
      (NMP_ComputeSoftmaxExp_for_asn_26_itm_2[25:0]), NMP_ComputeSoftmaxMax_for_if_less_4_itm);
  assign max_value_26_0_sva_dfm_10_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_9_1_26,
      (NMP_ComputeSoftmaxExp_for_asn_25_itm_2[26]), NMP_ComputeSoftmaxMax_for_if_less_5_itm_1);
  assign max_value_26_0_sva_dfm_10_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_9_1_25_0,
      (NMP_ComputeSoftmaxExp_for_asn_25_itm_2[25:0]), NMP_ComputeSoftmaxMax_for_if_less_5_itm_1);
  assign max_value_26_0_sva_dfm_8_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_7_26_mx0,
      (NMP_ComputeSoftmaxExp_for_asn_23_itm_1[26]), NMP_ComputeSoftmaxMax_for_if_less_7_itm);
  assign max_value_26_0_sva_dfm_8_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_7_25_0_mx0,
      (NMP_ComputeSoftmaxExp_for_asn_23_itm_1[25:0]), NMP_ComputeSoftmaxMax_for_if_less_7_itm);
  assign max_value_26_0_sva_dfm_7_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_6_1_26,
      (NMP_ComputeSoftmaxExp_for_asn_22_itm_1[26]), NMP_ComputeSoftmaxMax_for_if_less_8_itm);
  assign max_value_26_0_sva_dfm_7_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_6_1_25_0,
      (NMP_ComputeSoftmaxExp_for_asn_22_itm_1[25:0]), NMP_ComputeSoftmaxMax_for_if_less_8_itm);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_60_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_60_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_64_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_1_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_64_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_56_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_15_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_56_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_4_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_2_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_4_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_52_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_14_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_52_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_8_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_3_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_8_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_48_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_13_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_48_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_12_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_4_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_12_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_44_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_12_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_44_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_16_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_5_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_16_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_40_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_11_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_40_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_20_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_6_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_20_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_36_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_10_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_36_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_24_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_7_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_24_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_32_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_32_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z[31:22]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_28_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z[33:32]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_8_sva_1
      = ({ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_28_nl
      , 1'b0 , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z[32])
      , (~ (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z[33]))
      , (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z[33])})
      * (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z[31:22]);
  assign max_value_26_0_sva_dfm_5_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_4_26_mx0,
      (input_fixed_5_26_0_sva[26]), NMP_ComputeSoftmaxMax_for_if_less_10_itm);
  assign max_value_26_0_sva_dfm_5_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_4_25_0_mx0,
      (input_fixed_5_26_0_sva[25:0]), NMP_ComputeSoftmaxMax_for_if_less_10_itm);
  assign max_value_26_0_sva_dfm_4_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_3_26_mx0,
      (input_fixed_4_26_0_sva[26]), NMP_ComputeSoftmaxMax_for_if_less_11_itm);
  assign max_value_26_0_sva_dfm_4_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_3_25_0_mx0,
      (input_fixed_4_26_0_sva[25:0]), NMP_ComputeSoftmaxMax_for_if_less_11_itm);
  assign max_value_26_0_sva_dfm_3_26_mx0 = MUX_s_1_2_2(max_value_26_0_sva_dfm_2_1_26,
      (input_fixed_3_26_0_sva[26]), NMP_ComputeSoftmaxMax_for_if_less_12_itm_1);
  assign max_value_26_0_sva_dfm_3_25_0_mx0 = MUX_v_26_2_2(max_value_26_0_sva_dfm_2_1_25_0,
      (input_fixed_3_26_0_sva[25:0]), NMP_ComputeSoftmaxMax_for_if_less_12_itm_1);
  assign max_value_26_0_sva_dfm_1_26_1 = (input_fixed_1_26_0_sva[26]) & NMP_ComputeSoftmaxMax_for_if_less_14_ssc_1;
  assign max_value_26_0_sva_dfm_1_25_0_mx0 = MUX_v_26_2_2(NMP_ComputeSoftmaxMax_for_NMP_ComputeSoftmaxMax_for_and_psp_1,
      (input_fixed_1_26_0_sva[25:0]), NMP_ComputeSoftmaxMax_for_if_less_14_ssc_1);
  assign NMP_ComputeSoftmaxMax_for_if_less_14_ssc_1 = $signed({1'b0, NMP_ComputeSoftmaxMax_for_NMP_ComputeSoftmaxMax_for_and_psp_1})
      < $signed(input_fixed_1_26_0_sva);
  assign NMP_ComputeSoftmaxMax_for_NMP_ComputeSoftmaxMax_for_and_psp_1 = MUX_v_26_2_2(26'b00000000000000000000000000,
      (input_fixed_0_26_0_sva[25:0]), ($signed(1'b0) < $signed(input_fixed_0_26_0_sva)));
  assign nmp_config_ConfigRead_nor_2_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:1]!=15'b000000000000000));
  assign while_mux_1001_nl = MUX_s_1_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_54_itm,
      max_value_26_0_sva_26, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign max_value_mux_1_itm = MUX_s_1_2_2(max_value_26_0_sva_26, while_mux_1001_nl,
      while_stage_0_7);
  assign max_value_and_11_nl = (~ or_924_itm) & while_stage_0_7;
  assign max_value_mux_2_itm = MUX_v_26_2_2(max_value_26_0_sva_25_0, NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_52_itm,
      max_value_and_11_nl);
  assign while_asn_728 = NMP_RunFSM_switch_lp_equal_tmp_18 | NMP_RunFSM_switch_lp_equal_tmp_1_17
      | NMP_RunFSM_switch_lp_equal_tmp_2_17 | NMP_RunFSM_switch_lp_equal_tmp_3_17
      | NMP_RunFSM_switch_lp_equal_tmp_5_17 | NMP_RunFSM_switch_lp_equal_tmp_6_17
      | NMP_RunFSM_switch_lp_equal_tmp_7_17 | NMP_RunFSM_switch_lp_equal_tmp_9_17
      | NMP_RunFSM_switch_lp_equal_tmp_10_18 | NMP_RunFSM_switch_lp_equal_tmp_11_18
      | NMP_RunFSM_switch_lp_equal_tmp_12_18 | NMP_RunFSM_switch_lp_or_tmp_17 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_18;
  assign while_asn_730 = NMP_RunFSM_switch_lp_equal_tmp_4_17 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_18);
  assign while_asn_732 = NMP_RunFSM_switch_lp_equal_tmp_8_17 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_18);
  assign while_asn_734 = NMP_RunFSM_switch_lp_equal_tmp_17_1 | NMP_RunFSM_switch_lp_equal_tmp_1_16
      | NMP_RunFSM_switch_lp_equal_tmp_2_16 | NMP_RunFSM_switch_lp_equal_tmp_3_16
      | NMP_RunFSM_switch_lp_equal_tmp_5_16 | NMP_RunFSM_switch_lp_equal_tmp_6_16
      | NMP_RunFSM_switch_lp_equal_tmp_7_16 | NMP_RunFSM_switch_lp_equal_tmp_9_16
      | NMP_RunFSM_switch_lp_equal_tmp_10_17 | NMP_RunFSM_switch_lp_equal_tmp_11_17
      | NMP_RunFSM_switch_lp_equal_tmp_12_17 | NMP_RunFSM_switch_lp_or_tmp_16 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17;
  assign while_asn_736 = NMP_RunFSM_switch_lp_equal_tmp_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_asn_738 = NMP_RunFSM_switch_lp_equal_tmp_4_16 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17);
  assign while_asn_740 = NMP_RunFSM_switch_lp_equal_tmp_8_16 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17);
  assign out_adp_set_value_ac_float_mux_95_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_94_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_15_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_15_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_93_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_14_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_14_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_92_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_13_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_13_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_91_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_12_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_12_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_90_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_11_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_11_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_89_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_10_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_10_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_88_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_9_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_9_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_87_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_8_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_8_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_86_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_7_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_7_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_85_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_6_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_6_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_84_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_5_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_5_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_83_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_4_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_4_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_82_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_3_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_3_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_81_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_2_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_2_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_mux_80_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_ac_int_cctor_4_1_1_sva_1[3]),
      (out_adp_set_value_ac_float_exp_tmp_1_sva_2[4]), NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs);
  assign out_adp_set_value_ac_float_1_mux_95_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_94_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_15_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_15_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_93_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_14_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_14_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_92_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_13_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_13_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_91_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_12_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_12_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_90_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_11_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_11_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_89_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_10_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_10_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_88_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_9_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_9_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_87_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_8_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_8_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_86_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_7_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_7_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_85_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_6_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_6_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_84_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_5_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_5_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_83_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_4_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_4_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_82_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_3_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_3_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_81_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_2_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_2_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign out_adp_set_value_ac_float_1_mux_80_tmp_3 = MUX_s_1_2_2((out_adp_set_value_ac_float_1_ac_int_cctor_4_1_1_sva_1[3]),
      (out_adp_set_value_ac_float_1_exp_tmp_1_sva_2[4]), NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs);
  assign and_dcpl = while_stage_0_19 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17);
  assign and_dcpl_3 = NMP_RunFSM_switch_lp_conc_itm_16_0 & (~ NMP_RunFSM_switch_lp_conc_itm_16_2);
  assign and_dcpl_5 = while_stage_0_18 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_16);
  assign and_dcpl_6 = and_dcpl_5 & (~ NMP_RunFSM_switch_lp_conc_itm_16_1);
  assign and_dcpl_8 = NMP_RunFSM_switch_lp_conc_itm_16_2 & (~ NMP_RunFSM_switch_lp_conc_itm_16_3);
  assign and_dcpl_9 = (~ NMP_RunFSM_switch_lp_conc_itm_16_1) & NMP_RunFSM_switch_lp_conc_itm_16_0;
  assign and_dcpl_10 = and_dcpl_9 & and_dcpl_8;
  assign or_dcpl_5 = (NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_12 = (NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_19 = (NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_26 = (NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_33 = (NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_40 = (NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_47 = (NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_54 = (NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_61 = (NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_68 = (NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_75 = (NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_82 = (NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_89 = (NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_96 = (NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_103 = (NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_110 = (NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp!=7'b0000000);
  assign and_dcpl_46 = (~ NMP_RunFSM_switch_lp_conc_itm_16_2) & NMP_RunFSM_switch_lp_conc_itm_16_3;
  assign and_dcpl_47 = and_dcpl_9 & and_dcpl_46;
  assign or_dcpl_117 = (NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_124 = (NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_131 = (NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_138 = (NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_145 = (NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_152 = (NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_159 = (NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_166 = (NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_173 = (NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_180 = (NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_187 = (NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_194 = (NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_201 = (NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_208 = (NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_215 = (NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign or_dcpl_222 = (NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp!=7'b0000000);
  assign and_dcpl_88 = ~(NMP_RunFSM_switch_lp_conc_itm_15_1 | NMP_RunFSM_switch_lp_conc_itm_15_3);
  assign and_dcpl_90 = while_stage_0_17 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_15);
  assign and_dcpl_91 = and_dcpl_90 & NMP_RunFSM_switch_lp_conc_itm_15_0;
  assign and_dcpl_96 = while_stage_0_16 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_14);
  assign and_dcpl_97 = while_stage_0_15 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_13);
  assign and_dcpl_100 = while_stage_0_14 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_12);
  assign and_dcpl_101 = and_dcpl_100 & (~ NMP_RunFSM_switch_lp_conc_itm_12_1);
  assign and_dcpl_105 = NMP_RunFSM_switch_lp_conc_itm_12_3 & (~ NMP_RunFSM_switch_lp_conc_itm_12_2);
  assign and_dcpl_108 = and_dcpl_100 & (~ NMP_RunFSM_switch_lp_equal_tmp_12);
  assign and_dcpl_122 = NMP_RunFSM_switch_lp_conc_itm_11_2 & (~ NMP_RunFSM_switch_lp_conc_itm_11_3);
  assign and_dcpl_124 = while_stage_0_13 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11);
  assign and_dcpl_125 = and_dcpl_124 & (~ NMP_RunFSM_switch_lp_conc_itm_11_1);
  assign and_dcpl_129 = (~ NMP_RunFSM_switch_lp_conc_itm_11_2) & NMP_RunFSM_switch_lp_conc_itm_11_3;
  assign and_dcpl_130 = and_dcpl_129 & (~ NMP_RunFSM_switch_lp_conc_itm_11_0);
  assign and_dcpl_134 = ~(NMP_RunFSM_switch_lp_conc_itm_10_3 | NMP_RunFSM_switch_lp_conc_itm_10_1);
  assign and_dcpl_136 = while_stage_0_12 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10);
  assign and_dcpl_137 = and_dcpl_136 & NMP_RunFSM_switch_lp_conc_itm_10_2;
  assign and_dcpl_139 = NMP_RunFSM_switch_lp_conc_itm_10_3 & (~ NMP_RunFSM_switch_lp_conc_itm_10_1);
  assign and_dcpl_141 = and_dcpl_136 & (~ NMP_RunFSM_switch_lp_conc_itm_10_2);
  assign and_dcpl_142 = and_dcpl_141 & and_dcpl_139 & (~ NMP_RunFSM_switch_lp_conc_itm_10_0);
  assign and_dcpl_143 = ~(NMP_RunFSM_switch_lp_conc_itm_9_3 | NMP_RunFSM_switch_lp_conc_itm_9_1);
  assign and_dcpl_145 = while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9);
  assign and_dcpl_146 = and_dcpl_145 & NMP_RunFSM_switch_lp_conc_itm_9_2;
  assign and_dcpl_148 = NMP_RunFSM_switch_lp_conc_itm_9_3 & (~ NMP_RunFSM_switch_lp_conc_itm_9_1);
  assign and_dcpl_150 = and_dcpl_145 & (~ NMP_RunFSM_switch_lp_conc_itm_9_2);
  assign and_dcpl_152 = ~(NMP_RunFSM_switch_lp_conc_itm_8_1 | NMP_RunFSM_switch_lp_conc_itm_8_3);
  assign and_dcpl_154 = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign and_dcpl_155 = and_dcpl_154 & NMP_RunFSM_switch_lp_conc_itm_8_2;
  assign and_dcpl_159 = while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign and_dcpl_162 = while_stage_0_8 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6);
  assign and_dcpl_163 = while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_dcpl_164 = NMP_RunFSM_switch_lp_conc_itm_4_2 & NMP_RunFSM_switch_lp_conc_itm_4_1;
  assign and_dcpl_166 = while_stage_0_6 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_dcpl_167 = and_dcpl_166 & (~ NMP_RunFSM_switch_lp_conc_itm_4_3);
  assign and_dcpl_169 = while_stage_0_5 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_3);
  assign and_dcpl_170 = while_stage_0_4 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign and_dcpl_171 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign or_tmp = state_2_sva | state_0_sva;
  assign and_dcpl_172 = reg_rva_in_PopNB_mioi_iswt0_cse & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign or_tmp_12 = NMP_UpdateFSM_switch_lp_equal_tmp_5_1 | NMP_UpdateFSM_switch_lp_equal_tmp_6_1;
  assign nand_3_nl = ~(state_1_sva & state_3_sva & (~ state_2_sva) & state_0_sva);
  assign nor_45_nl = ~(NMP_UpdateFSM_switch_lp_equal_tmp_3_1 | NMP_UpdateFSM_switch_lp_equal_tmp_2_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_1_1 | (~(or_tmp_12 | (~(NMP_UpdateFSM_switch_lp_or_tmp_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_4_1 | NMP_UpdateFSM_switch_lp_equal_tmp_1
      | NMP_UpdateFSM_switch_lp_nor_tmp_1 | NMP_RunFSM_switch_lp_equal_tmp_12_1 |
      NMP_RunFSM_switch_lp_equal_tmp_1 | NMP_RunFSM_switch_lp_equal_tmp_11_1 | (~
      next_state_3_lpi_1_dfm_3) | (~ NMP_RunFSM_switch_lp_or_73_tmp) | (~ state_0_sva)
      | state_2_sva)))));
  assign nor_46_nl = ~((~ state_3_sva) | state_2_sva | (~ state_0_sva));
  assign mux_5_nl = MUX_s_1_2_2(nor_45_nl, nor_46_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nand_nl = ~(state_1_sva_dfm_1 & mux_5_nl);
  assign mux_tmp_6 = MUX_s_1_2_2(nand_3_nl, nand_nl, while_stage_0_3);
  assign and_dcpl_176 = and_dcpl_5 & and_dcpl_9;
  assign and_dcpl_177 = and_dcpl_176 & and_dcpl_8 & NMP_RunFSM_switch_lp_equal_tmp_4_15;
  assign and_dcpl_195 = and_dcpl_176 & and_dcpl_46 & NMP_RunFSM_switch_lp_equal_tmp_8_15;
  assign and_dcpl_213 = NMP_RunFSM_switch_lp_conc_itm_15_0 & (~ NMP_RunFSM_switch_lp_conc_itm_15_1);
  assign or_dcpl_309 = (and_dcpl_213 & (~(NMP_RunFSM_switch_lp_conc_itm_15_3 | NMP_RunFSM_switch_lp_conc_itm_15_2)))
      | (~(NMP_RunFSM_switch_lp_equal_tmp_9_14 & while_stage_0_17)) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_15;
  assign and_dcpl_215 = (~ NMP_RunFSM_switch_lp_conc_itm_15_3) & NMP_RunFSM_switch_lp_conc_itm_15_2;
  assign and_dcpl_217 = and_dcpl_90 & and_dcpl_213;
  assign and_dcpl_249 = NMP_RunFSM_switch_lp_conc_itm_15_3 & (~ NMP_RunFSM_switch_lp_conc_itm_15_2);
  assign and_dcpl_283 = and_dcpl_159 & (~ NMP_RunFSM_switch_lp_conc_itm_7_3) & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign or_tmp_21 = (~ NMP_RunFSM_switch_lp_conc_itm_7_1) | NMP_RunFSM_switch_lp_equal_tmp_7
      | (~ NMP_RunFSM_switch_lp_equal_tmp_6_6);
  assign mux_tmp_7 = MUX_s_1_2_2(NMP_RunFSM_switch_lp_conc_itm_7_1, or_tmp_21, NMP_RunFSM_switch_lp_conc_itm_7_0);
  assign and_dcpl_292 = and_dcpl_167 & and_dcpl_164 & (~ NMP_RunFSM_switch_lp_conc_itm_4_0);
  assign and_dcpl_293 = NMP_RunFSM_switch_lp_conc_itm_3_2 & NMP_RunFSM_switch_lp_conc_itm_3_1;
  assign and_dcpl_295 = and_dcpl_169 & (~ NMP_RunFSM_switch_lp_conc_itm_3_3);
  assign and_dcpl_296 = and_dcpl_295 & and_dcpl_293 & NMP_RunFSM_switch_lp_conc_itm_3_0;
  assign and_dcpl_298 = (~ NMP_RunFSM_switch_lp_conc_itm_8_1) & NMP_RunFSM_switch_lp_conc_itm_8_3;
  assign and_dcpl_300 = and_dcpl_154 & (~ NMP_RunFSM_switch_lp_conc_itm_8_2);
  assign and_dcpl_305 = and_dcpl_162 & (~ NMP_RunFSM_switch_lp_conc_itm_6_1);
  assign and_dcpl_317 = and_dcpl_124 & (~ NMP_RunFSM_switch_lp_equal_tmp_11);
  assign and_dcpl_320 = and_dcpl_134 & NMP_RunFSM_switch_lp_conc_itm_10_0;
  assign and_dcpl_342 = and_dcpl_295 & and_dcpl_293 & (~ NMP_RunFSM_switch_lp_conc_itm_3_0);
  assign and_dcpl_343 = NMP_RunFSM_switch_lp_conc_itm_3_1 & (~ NMP_RunFSM_switch_lp_conc_itm_3_0);
  assign and_dcpl_346 = and_dcpl_169 & (~ NMP_RunFSM_switch_lp_conc_itm_3_3) & NMP_RunFSM_switch_lp_conc_itm_3_2;
  assign and_dcpl_354 = and_dcpl_163 & (~ NMP_RunFSM_switch_lp_conc_itm_5_1);
  assign and_dcpl_360 = NMP_RunFSM_switch_lp_conc_itm_14_0 & (~ NMP_RunFSM_switch_lp_conc_itm_14_2);
  assign and_dcpl_362 = and_dcpl_96 & (~ NMP_RunFSM_switch_lp_conc_itm_14_1);
  assign and_dcpl_365 = and_dcpl_150 & and_dcpl_148 & NMP_RunFSM_switch_lp_conc_itm_9_0;
  assign and_dcpl_367 = and_dcpl_170 & (~ NMP_RunFSM_switch_lp_conc_itm_2_3);
  assign and_dcpl_369 = NMP_RunFSM_switch_lp_conc_itm_2_2 & NMP_RunFSM_switch_lp_conc_itm_2_0;
  assign and_dcpl_376 = and_dcpl_143 & NMP_RunFSM_switch_lp_conc_itm_9_0;
  assign and_dcpl_377 = and_dcpl_146 & and_dcpl_376;
  assign and_dcpl_409 = NMP_RunFSM_switch_lp_conc_itm_4_2 & (~ NMP_RunFSM_switch_lp_conc_itm_4_1);
  assign and_dcpl_418 = and_dcpl_97 & (~ NMP_RunFSM_switch_lp_conc_itm_13_1);
  assign and_dcpl_424 = NMP_RunFSM_switch_lp_conc_itm_13_0 & (~ NMP_RunFSM_switch_lp_conc_itm_13_3);
  assign and_dcpl_427 = and_dcpl_152 & NMP_RunFSM_switch_lp_conc_itm_8_0;
  assign and_dcpl_440 = NMP_RunFSM_switch_lp_conc_itm_3_2 & (~ NMP_RunFSM_switch_lp_conc_itm_3_1);
  assign and_dcpl_443 = state_1_sva & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign and_dcpl_482 = NMP_RunFSM_switch_lp_conc_itm_5_0 & (~ NMP_RunFSM_switch_lp_conc_itm_5_3);
  assign and_dcpl_492 = and_dcpl_167 & and_dcpl_409 & NMP_RunFSM_switch_lp_conc_itm_4_0;
  assign and_dcpl_504 = and_dcpl_295 & and_dcpl_440 & NMP_RunFSM_switch_lp_conc_itm_3_0;
  assign and_dcpl_509 = and_dcpl_367 & and_dcpl_369 & (~ NMP_RunFSM_switch_lp_conc_itm_2_1);
  assign and_dcpl_519 = NMP_RunFSM_switch_lp_conc_itm_6_0 & (~ NMP_RunFSM_switch_lp_conc_itm_6_2);
  assign and_dcpl_541 = and_dcpl_166 & NMP_RunFSM_switch_lp_conc_itm_4_3;
  assign and_dcpl_544 = (~(NMP_RunFSM_switch_lp_conc_itm_4_2 | NMP_RunFSM_switch_lp_conc_itm_4_1))
      & NMP_RunFSM_switch_lp_conc_itm_4_0;
  assign and_dcpl_554 = and_dcpl_169 & NMP_RunFSM_switch_lp_conc_itm_3_3;
  assign and_dcpl_557 = (~(NMP_RunFSM_switch_lp_conc_itm_3_2 | NMP_RunFSM_switch_lp_conc_itm_3_1))
      & NMP_RunFSM_switch_lp_conc_itm_3_0;
  assign and_dcpl_564 = and_dcpl_170 & NMP_RunFSM_switch_lp_conc_itm_2_3;
  assign and_dcpl_567 = (~ NMP_RunFSM_switch_lp_conc_itm_2_2) & NMP_RunFSM_switch_lp_conc_itm_2_0
      & (~ NMP_RunFSM_switch_lp_conc_itm_2_1);
  assign and_dcpl_581 = fsm_output & (~ NMP_RunFSM_switch_lp_conc_itm_17_0);
  assign or_tmp_35 = (~ NMP_RunFSM_switch_lp_conc_itm_2_1) | (~ NMP_RunFSM_switch_lp_conc_itm_2_0)
      | NMP_RunFSM_switch_lp_conc_itm_2_2 | NMP_RunFSM_switch_lp_conc_itm_2_3 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4);
  assign or_tmp_40 = NMP_RunFSM_switch_lp_conc_itm_14_3 | (~ NMP_RunFSM_switch_lp_conc_itm_14_2)
      | (~ NMP_RunFSM_switch_lp_conc_itm_14_0) | NMP_RunFSM_switch_lp_conc_itm_14_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_14
      | (~ while_stage_0_16);
  assign nor_79_nl = ~(while_stage_0_15 | (~ or_tmp_40));
  assign or_509_nl = (~ NMP_RunFSM_switch_lp_conc_itm_13_2) | NMP_RunFSM_switch_lp_conc_itm_13_3
      | (~ NMP_RunFSM_switch_lp_conc_itm_13_0) | NMP_RunFSM_switch_lp_conc_itm_13_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_13;
  assign mux_tmp_17 = MUX_s_1_2_2(nor_79_nl, or_tmp_40, or_509_nl);
  assign or_tmp_45 = (~ NMP_RunFSM_switch_lp_conc_itm_5_2) | NMP_RunFSM_switch_lp_conc_itm_5_3
      | (~ NMP_RunFSM_switch_lp_conc_itm_5_0) | (~ NMP_RunFSM_switch_lp_conc_itm_5_1)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7);
  assign or_tmp_50 = (~ NMP_RunFSM_switch_lp_conc_itm_14_3) | NMP_RunFSM_switch_lp_conc_itm_14_2
      | (~ NMP_RunFSM_switch_lp_conc_itm_14_0) | NMP_RunFSM_switch_lp_conc_itm_14_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_14
      | (~ while_stage_0_16);
  assign nor_80_nl = ~(while_stage_0_15 | (~ or_tmp_50));
  assign or_519_nl = NMP_RunFSM_switch_lp_conc_itm_13_2 | (~ NMP_RunFSM_switch_lp_conc_itm_13_3)
      | (~ NMP_RunFSM_switch_lp_conc_itm_13_0) | NMP_RunFSM_switch_lp_conc_itm_13_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_13;
  assign mux_tmp_20 = MUX_s_1_2_2(nor_80_nl, or_tmp_50, or_519_nl);
  assign or_tmp_56 = (state_0_sva & NMP_RunFSM_switch_lp_or_73_tmp) | NMP_RunFSM_switch_lp_equal_tmp_12_1;
  assign or_tmp_57 = (~ or_tmp_56) | NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign or_tmp_60 = (~((or_tmp & NMP_RunFSM_switch_lp_or_73_tmp) | NMP_RunFSM_switch_lp_equal_tmp_12_1))
      | NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign mux_280_nl = MUX_s_1_2_2(or_tmp_60, or_803_cse, next_state_3_lpi_1_dfm_3);
  assign mux_tmp_25 = MUX_s_1_2_2(mux_280_nl, or_tmp_60, NMP_RunFSM_switch_lp_equal_tmp_11_1);
  assign mux_tmp_26 = MUX_s_1_2_2(mux_tmp_25, or_tmp_57, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign or_tmp_85 = state_2_sva | state_1_sva | state_0_sva | state_3_sva;
  assign or_tmp_87 = NMP_RunFSM_switch_lp_conc_itm_17_1 | (~ NMP_RunFSM_switch_lp_conc_itm_17_0);
  assign or_dcpl_471 = (~ while_stage_0_19) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17;
  assign or_dcpl_475 = (~(rva_in_PopNB_mioi_return_rsc_z_mxwt & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt))
      | nmp_config_ConfigRead_unequal_tmp_1;
  assign or_dcpl_477 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]));
  assign or_dcpl_480 = or_dcpl_477 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) & reg_rva_in_PopNB_mioi_iswt0_cse))
      | or_dcpl_475;
  assign or_dcpl_481 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ while_stage_0_3);
  assign or_dcpl_483 = NMP_RunFSM_switch_lp_conc_itm_17_3 | (~ NMP_RunFSM_switch_lp_conc_itm_17_2);
  assign or_dcpl_485 = or_dcpl_471 | or_tmp_87;
  assign or_dcpl_489 = or_tmp_87 | NMP_RunFSM_switch_lp_conc_itm_17_3;
  assign or_dcpl_582 = (~ NMP_RunFSM_switch_lp_conc_itm_17_3) | NMP_RunFSM_switch_lp_conc_itm_17_2;
  assign or_dcpl_587 = or_tmp_87 | (~ NMP_RunFSM_switch_lp_conc_itm_17_3);
  assign or_dcpl_679 = (~ while_stage_0_18) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_16;
  assign or_dcpl_684 = (~ while_stage_0_14) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_12
      | NMP_RunFSM_switch_lp_conc_itm_12_1;
  assign and_dcpl_634 = (ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_3==40'b0000000000000000000000000000000000000000);
  assign NMP_ComputeSoftmaxMax_for_if_less_2_itm = $signed(({max_value_26_0_sva_dfm_12_26_mx0
      , max_value_26_0_sva_dfm_12_25_0_mx0})) < $signed(NMP_ComputeSoftmaxExp_for_asn_28_itm_2);
  assign or_dcpl_694 = or_dcpl_477 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]));
  assign or_tmp_89 = (~ state_0_sva) | state_1_sva_dfm_1;
  assign or_tmp_90 = state_0_sva | (~ state_1_sva_dfm_1);
  assign or_tmp_91 = NMP_UpdateFSM_switch_lp_equal_tmp_4_1 | NMP_UpdateFSM_switch_lp_or_tmp_1;
  assign or_tmp_92 = NMP_UpdateFSM_switch_lp_equal_tmp_2_1 | NMP_UpdateFSM_switch_lp_equal_tmp_3_1
      | state_1_sva_dfm_1;
  assign or_tmp_95 = NMP_UpdateFSM_switch_lp_equal_tmp_2_1 | NMP_UpdateFSM_switch_lp_equal_tmp_3_1;
  assign or_tmp_96 = state_1_sva_dfm_1 | NMP_UpdateFSM_switch_lp_equal_tmp_5_1 |
      NMP_UpdateFSM_switch_lp_equal_tmp_6_1;
  assign mux_tmp_83 = MUX_s_1_2_2((~ or_tmp_12), or_tmp_12, state_1_sva_dfm_1);
  assign or_tmp_99 = state_1_sva_dfm_1 | (~ or_tmp_12);
  assign mux_tmp_85 = MUX_s_1_2_2(state_1_sva_dfm_1, mux_tmp_83, or_803_cse);
  assign or_799_nl = (~ state_2_sva) | (~ NMP_RunFSM_switch_lp_or_73_tmp) | NMP_UpdateFSM_switch_lp_equal_tmp_1
      | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign mux_tmp_89 = MUX_s_1_2_2(state_1_sva_dfm_1, mux_tmp_83, or_799_nl);
  assign nor_16_nl = ~(state_2_sva | (~ NMP_RunFSM_switch_lp_or_73_tmp));
  assign mux_98_nl = MUX_s_1_2_2(mux_110_cse, mux_tmp_85, nor_16_nl);
  assign mux_tmp_99 = MUX_s_1_2_2(mux_tmp_89, mux_98_nl, next_state_3_lpi_1_dfm_3);
  assign nor_tmp_17 = state_0_sva & state_1_sva;
  assign or_tmp_116 = (~ NMP_RunFSM_switch_lp_equal_tmp_11_1) | NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2;
  assign mux_tmp_139 = MUX_s_1_2_2(or_tmp_89, or_tmp_90, state_3_sva);
  assign or_819_nl = (~ state_0_sva) | state_1_sva;
  assign or_818_nl = state_0_sva | (~ state_1_sva);
  assign mux_tmp_140 = MUX_s_1_2_2(or_819_nl, or_818_nl, state_3_sva);
  assign nor_tmp_19 = or_tmp_91 & state_1_sva_dfm_1;
  assign mux_tmp_142 = MUX_s_1_2_2((~ state_1_sva_dfm_1), state_1_sva_dfm_1, or_tmp_91);
  assign or_823_nl = (~(NMP_RunFSM_switch_lp_equal_tmp_12_1 | NMP_RunFSM_switch_lp_or_73_tmp))
      | NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign mux_tmp_143 = MUX_s_1_2_2(mux_tmp_142, nor_tmp_19, or_823_nl);
  assign or_tmp_129 = and_899_cse | NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign or_827_nl = state_2_sva | (~ NMP_RunFSM_switch_lp_or_73_tmp) | NMP_UpdateFSM_switch_lp_equal_tmp_1
      | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign mux_tmp_147 = MUX_s_1_2_2(mux_tmp_142, nor_tmp_19, or_827_nl);
  assign mux_tmp_150 = MUX_s_1_2_2(mux_149_itm, mux_tmp_147, NMP_RunFSM_switch_lp_equal_tmp_11_1);
  assign mux_tmp_151 = MUX_s_1_2_2(mux_tmp_150, mux_219_cse, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign mux_tmp_152 = MUX_s_1_2_2(mux_tmp_151, mux_tmp_143, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_tmp_156 = MUX_s_1_2_2(mux_tmp_142, nor_tmp_19, or_533_cse);
  assign mux_tmp_161 = MUX_s_1_2_2(mux_tmp_142, nor_tmp_19, or_803_cse);
  assign not_tmp_277 = ~(state_0_sva | (~ reg_rva_in_PopNB_mioi_iswt0_cse));
  assign or_tmp_147 = state_1_sva_dfm_1 | (~ reg_rva_in_PopNB_mioi_iswt0_cse);
  assign nor_tmp_31 = or_tmp_85 & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign not_tmp_279 = ~(state_0_sva & reg_rva_in_PopNB_mioi_iswt0_cse);
  assign or_tmp_159 = nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1
      | operator_16_false_acc_2_itm_17 | (~ state_1_sva) | (~ state_3_sva) | state_2_sva
      | not_tmp_279;
  assign or_tmp_165 = (~ large_rsp_PopNB_mioi_return_rsc_z_mxwt) | (~ state_1_sva)
      | state_3_sva | state_2_sva | state_0_sva;
  assign not_tmp_286 = ~(or_tmp_165 | (~ reg_rva_in_PopNB_mioi_iswt0_cse));
  assign or_dcpl_700 = or_dcpl_679 | NMP_RunFSM_switch_lp_conc_itm_16_1;
  assign or_dcpl_708 = (~ while_stage_0_13) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11
      | NMP_RunFSM_switch_lp_conc_itm_11_1;
  assign NMP_ComputeSoftmaxMax_for_if_less_6_itm = $signed(({max_value_26_0_sva_dfm_8_26_mx0
      , max_value_26_0_sva_dfm_8_25_0_mx0})) < $signed(NMP_ComputeSoftmaxExp_for_asn_24_itm_1);
  assign and_dcpl_750 = (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]);
  assign or_dcpl_718 = (~ while_stage_0_12) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10;
  assign and_dcpl_832 = ~(NMP_RunFSM_switch_lp_conc_itm_7_3 | NMP_RunFSM_switch_lp_conc_itm_7_1);
  assign NMP_ComputeSoftmaxMax_for_if_less_9_itm = $signed(({max_value_26_0_sva_dfm_5_26_mx0
      , max_value_26_0_sva_dfm_5_25_0_mx0})) < $signed(input_fixed_6_26_0_sva);
  assign NMP_ComputeSoftmaxMax_for_if_less_13_itm = $signed(({max_value_26_0_sva_dfm_1_26_1
      , max_value_26_0_sva_dfm_1_25_0_mx0})) < $signed(input_fixed_2_26_0_sva);
  assign NMP_ComputeSoftmaxMax_for_if_less_1_itm = $signed(({max_value_26_0_sva_dfm_13_1_26
      , max_value_26_0_sva_dfm_13_1_25_0})) < $signed(NMP_ComputeSoftmaxMax_for_asn_13_itm_3);
  assign NMP_ComputeSoftmaxMax_for_if_less_3_itm = $signed(({max_value_26_0_sva_dfm_11_26_mx0
      , max_value_26_0_sva_dfm_11_25_0_mx0})) < $signed(NMP_ComputeSoftmaxExp_for_asn_27_itm_2);
  assign NMP_ComputeSoftmaxMax_for_if_less_4_itm = $signed(({max_value_26_0_sva_dfm_10_26_mx0
      , max_value_26_0_sva_dfm_10_25_0_mx0})) < $signed(NMP_ComputeSoftmaxExp_for_asn_26_itm_2);
  assign NMP_ComputeSoftmaxMax_for_if_less_7_itm = $signed(({max_value_26_0_sva_dfm_7_26_mx0
      , max_value_26_0_sva_dfm_7_25_0_mx0})) < $signed(NMP_ComputeSoftmaxExp_for_asn_23_itm_1);
  assign NMP_ComputeSoftmaxMax_for_if_less_8_itm = $signed(({max_value_26_0_sva_dfm_6_1_26
      , max_value_26_0_sva_dfm_6_1_25_0})) < $signed(NMP_ComputeSoftmaxExp_for_asn_22_itm_1);
  assign NMP_ComputeSoftmaxMax_for_if_less_10_itm = $signed(({max_value_26_0_sva_dfm_4_26_mx0
      , max_value_26_0_sva_dfm_4_25_0_mx0})) < $signed(input_fixed_5_26_0_sva);
  assign NMP_ComputeSoftmaxMax_for_if_less_11_itm = $signed(({max_value_26_0_sva_dfm_3_26_mx0
      , max_value_26_0_sva_dfm_3_25_0_mx0})) < $signed(input_fixed_4_26_0_sva);
  assign and_dcpl_875 = and_dcpl_750 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]);
  assign nmp_config_adpbias_1_sva_dfm_3_1_mx0c0 = and_dcpl_750 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) & reg_rva_in_PopNB_mioi_iswt0_cse
      & rva_in_PopNB_mioi_return_rsc_z_mxwt & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & nmp_config_ConfigRead_nor_2_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]);
  assign nmp_config_adpbias_1_sva_dfm_3_1_mx0c1 = (or_dcpl_694 | or_dcpl_475) & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign nmp_config_adpbias_1_sva_dfm_3_1_mx0c2 = (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      & while_stage_0_3;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_a = NMP_ComputeSoftmaxNormalize_for_asn_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_pff = sum_exp_reciprocal_mux_rmff;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_a = NMP_ComputeSoftmaxNormalize_for_asn_45_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_a = NMP_ComputeSoftmaxNormalize_for_asn_43_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_a = NMP_ComputeSoftmaxNormalize_for_asn_41_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_a = NMP_ComputeSoftmaxNormalize_for_asn_39_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_a = NMP_ComputeSoftmaxNormalize_for_asn_37_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_a = NMP_ComputeSoftmaxNormalize_for_asn_35_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_a = NMP_ComputeSoftmaxNormalize_for_asn_33_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_a = NMP_ComputeSoftmaxNormalize_for_asn_31_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_a = NMP_ComputeSoftmaxNormalize_for_asn_29_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_a = NMP_ComputeSoftmaxNormalize_for_asn_27_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_a = NMP_ComputeSoftmaxNormalize_for_asn_25_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_a = NMP_ComputeSoftmaxNormalize_for_asn_23_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_a = NMP_ComputeSoftmaxNormalize_for_asn_21_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_a = NMP_ComputeSoftmaxNormalize_for_asn_19_itm_4;
  assign NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_a = NMP_ComputeSoftmaxNormalize_for_asn_17_itm_4;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_b
      = NMP_ComputeSoftmaxExp_for_1_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_b
      = NMP_ComputeSoftmaxExp_for_16_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_b
      = NMP_ComputeSoftmaxExp_for_15_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_b
      = NMP_ComputeSoftmaxExp_for_14_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_b
      = NMP_ComputeSoftmaxExp_for_13_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_b
      = NMP_ComputeSoftmaxExp_for_12_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_b
      = NMP_ComputeSoftmaxExp_for_11_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_b
      = NMP_ComputeSoftmaxExp_for_10_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_b
      = NMP_ComputeSoftmaxExp_for_9_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_b
      = NMP_ComputeSoftmaxExp_for_8_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_b
      = NMP_ComputeSoftmaxExp_for_7_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_b
      = NMP_ComputeSoftmaxExp_for_6_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_b
      = NMP_ComputeSoftmaxExp_for_5_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_b
      = NMP_ComputeSoftmaxExp_for_4_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_b
      = NMP_ComputeSoftmaxExp_for_3_acc_1_itm_1;
  assign NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_b
      = NMP_ComputeSoftmaxExp_for_2_acc_1_itm_1;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_a = NMP_ComputeRMSNormalize_for_asn_itm_11;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_b_pff = rms_reciprocal_mux_rmff;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_1_a = NMP_ComputeRMSNormalize_for_asn_60_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_2_a = NMP_ComputeRMSNormalize_for_asn_58_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_3_a = NMP_ComputeRMSNormalize_for_asn_56_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_4_a = NMP_ComputeRMSNormalize_for_asn_54_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_5_a = NMP_ComputeRMSNormalize_for_asn_52_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_6_a = NMP_ComputeRMSNormalize_for_asn_50_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_7_a = NMP_ComputeRMSNormalize_for_asn_48_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_8_a = NMP_ComputeRMSNormalize_for_asn_46_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_9_a = NMP_ComputeRMSNormalize_for_asn_44_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_10_a = NMP_ComputeRMSNormalize_for_asn_42_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_11_a = NMP_ComputeRMSNormalize_for_asn_40_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_12_a = NMP_ComputeRMSNormalize_for_asn_38_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_13_a = NMP_ComputeRMSNormalize_for_asn_36_itm_10;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_14_a = NMP_ComputeRMSNormalize_for_asn_34_itm_11;
  assign NMP_ComputeRMSNormalize_for_1_mul_cmp_15_a = NMP_ComputeRMSNormalize_for_asn_32_itm_11;
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_a_pff = input_fixed_0_26_0_sva;
  assign input_fixed_and_37_cse = (~ while_stage_0_4) & fsm_output;
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_a_pff = MUX_v_27_2_2(input_fixed_11_26_0_sva_dfm_2_1,
      input_fixed_11_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_a_pff = MUX_v_27_2_2(input_fixed_10_26_0_sva_dfm_2_1,
      input_fixed_10_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_a_pff = MUX_v_27_2_2(input_fixed_9_26_0_sva_dfm_2_1,
      input_fixed_9_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_a_pff = MUX_v_27_2_2(input_fixed_8_26_0_sva_dfm_2_1,
      input_fixed_8_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_a_pff = MUX_v_27_2_2(input_fixed_7_26_0_sva_dfm_2_1,
      input_fixed_7_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_a_pff = MUX_v_27_2_2(input_fixed_6_26_0_sva_dfm_2_1,
      input_fixed_6_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_a_pff = MUX_v_27_2_2(input_fixed_5_26_0_sva_dfm_2_1,
      input_fixed_5_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_a_pff = MUX_v_27_2_2(input_fixed_4_26_0_sva_dfm_2_1,
      input_fixed_4_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_a_pff = MUX_v_27_2_2(input_fixed_3_26_0_sva_dfm_2_1,
      input_fixed_3_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_a_pff = MUX_v_27_2_2(input_fixed_15_26_0_sva_dfm_2_1,
      input_fixed_15_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_a_pff = MUX_v_27_2_2(input_fixed_14_26_0_sva_dfm_2_1,
      input_fixed_14_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_a_pff = MUX_v_27_2_2(input_fixed_13_26_0_sva_dfm_2_1,
      input_fixed_13_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_a_pff = MUX_v_27_2_2(input_fixed_12_26_0_sva_dfm_2_1,
      input_fixed_12_26_0_sva, input_fixed_and_37_cse);
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_a_pff = input_fixed_2_26_0_sva;
  assign NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_a_pff = input_fixed_1_26_0_sva;
  assign or_dcpl_742 = (~(NMP_RunFSM_switch_lp_equal_tmp_8 | NMP_RunFSM_switch_lp_equal_tmp_6_7))
      | (~ while_stage_0_10) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  assign and_dcpl_887 = fsm_output & NMP_RunFSM_switch_lp_conc_itm_11_3;
  assign and_dcpl_893 = (~ NMP_RunFSM_switch_lp_conc_itm_10_2) & fsm_output;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_enex5
      = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_2_cse
      & (reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo
      | reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_1
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo);
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_3_enex5
      = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_2_cse
      & (reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_1
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_1
      | reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_2
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_1);
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_4_enex5
      = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_2_cse
      & (reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_2
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_2
      | reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_3
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_2);
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_5_enex5
      = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_2_cse
      & (reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_3
      | reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_4
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_3
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_3);
  assign nand_5_nl = ~(NMP_RunFSM_switch_lp_conc_itm_7_0 & NMP_RunFSM_switch_lp_conc_itm_7_1
      & (~ NMP_RunFSM_switch_lp_equal_tmp_7) & NMP_RunFSM_switch_lp_equal_tmp_6_6);
  assign nor_1_nl = ~(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_0_3_itm_3
      | (~ (ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_3[0])));
  assign mux_8_nl = MUX_s_1_2_2(mux_tmp_7, nand_5_nl, nor_1_nl);
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc
      = NMPRun_wen & (~ mux_8_nl) & and_dcpl_283;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5
      = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc
      & (reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mux_1_itm_2_enexo
      | reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1_enexo);
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5
      = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc
      & reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1_enexo_1;
  assign or_452_nl = NMP_RunFSM_switch_lp_conc_itm_7_3 | NMP_RunFSM_switch_lp_equal_tmp_7
      | (~ NMP_RunFSM_switch_lp_equal_tmp_6_6);
  assign mux_9_nl = MUX_s_1_2_2(NMP_RunFSM_switch_lp_conc_itm_7_3, or_452_nl, NMP_RunFSM_switch_lp_conc_itm_7_1);
  assign mux_10_nl = MUX_s_1_2_2(NMP_RunFSM_switch_lp_conc_itm_7_1, mux_9_nl, NMP_RunFSM_switch_lp_conc_itm_7_2);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_29_ssc
      = NMPRun_wen & (~ mux_10_nl) & and_dcpl_159 & NMP_RunFSM_switch_lp_conc_itm_7_0;
  assign nor_54_nl = ~(NMP_RunFSM_switch_lp_conc_itm_7_2 | (~ NMP_RunFSM_switch_lp_conc_itm_7_3));
  assign nor_55_nl = ~((~ NMP_RunFSM_switch_lp_conc_itm_7_2) | NMP_RunFSM_switch_lp_conc_itm_7_3
      | NMP_RunFSM_switch_lp_equal_tmp_7 | (~ NMP_RunFSM_switch_lp_equal_tmp_6_6));
  assign mux_11_nl = MUX_s_1_2_2(nor_54_nl, nor_55_nl, NMP_RunFSM_switch_lp_conc_itm_7_0);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_36_ssc
      = NMPRun_wen & mux_11_nl & and_dcpl_159 & NMP_RunFSM_switch_lp_conc_itm_7_1;
  assign nor_58_cse = ~(NMP_RunFSM_switch_lp_conc_itm_5_1 | NMP_RunFSM_switch_lp_conc_itm_5_3);
  assign mux_12_nl = MUX_s_1_2_2(NMP_RunFSM_switch_lp_conc_itm_5_0, (~ NMP_RunFSM_switch_lp_conc_itm_5_0),
      NMP_RunFSM_switch_lp_conc_itm_5_2);
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc
      = NMPRun_wen & mux_12_nl & and_dcpl_163 & nor_58_cse;
  assign NMP_PrepareReadReq_and_63_enex5 = NMP_PrepareReadReq_and_23_cse & reg_NMP_PrepareReadReq_asn_1_itm_12_1_enexo;
  assign NMP_ComputeRMSSqrtRecip_variance_and_enex5 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_9_cse
      & reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_enexo;
  assign NMP_ComputeRMSSqrtRecip_variance_and_2_enex5 = ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_9_cse
      & reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_1_enexo_1;
  assign NMP_ComputeRMSSqrtRecip_variance_and_1_ssc = NMPRun_wen & and_dcpl_295 &
      and_dcpl_440;
  assign NMP_PrepareReadReq_and_64_enex5 = NMP_PrepareReadReq_and_26_cse & reg_NMP_PrepareReadReq_asn_1_itm_11_1_enexo;
  assign NMP_PrepareReadReq_and_65_enex5 = NMP_PrepareReadReq_and_29_ssc & reg_NMP_PrepareReadReq_asn_1_itm_10_1_enexo;
  assign NMP_PrepareWriteReq_and_78_enex5 = NMP_PrepareWriteReq_and_35_cse & reg_NMP_PrepareWriteReq_asn_2_itm_8_enexo;
  assign NMP_PrepareWriteReq_and_79_enex5 = NMP_PrepareWriteReq_and_35_cse & reg_NMP_PrepareWriteReq_asn_2_itm_8_1_enexo;
  assign out_adp_set_value_ac_float_1_and_7_ssc = NMPRun_wen & (and_dcpl_365 | and_dcpl_377);
  assign NMP_PrepareReadReq_and_66_enex5 = NMP_PrepareReadReq_and_36_cse & reg_NMP_PrepareReadReq_asn_2_itm_8_1_enexo;
  assign NMP_PrepareWriteReq_and_80_enex5 = NMP_PrepareWriteReq_and_38_cse & reg_NMP_PrepareWriteReq_asn_2_itm_7_enexo;
  assign NMP_PrepareWriteReq_and_81_enex5 = NMP_PrepareWriteReq_and_38_cse & reg_NMP_PrepareWriteReq_asn_2_itm_7_1_enexo;
  assign out_adp_set_value_ac_float_1_and_8_ssc = NMPRun_wen & (NMP_RunFSM_switch_lp_conc_itm_8_2
      ^ NMP_RunFSM_switch_lp_conc_itm_8_3) & while_stage_0_10 & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
      | NMP_RunFSM_switch_lp_conc_itm_8_1)) & NMP_RunFSM_switch_lp_conc_itm_8_0;
  assign NMP_PrepareReadReq_and_67_enex5 = NMP_PrepareReadReq_and_39_cse & reg_NMP_PrepareReadReq_asn_2_itm_7_1_enexo;
  assign NMP_PrepareWriteReq_and_82_enex5 = ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_36_ssc
      & reg_NMP_PrepareWriteReq_asn_2_itm_6_enexo;
  assign mux_13_nl = MUX_s_1_2_2(NMP_RunFSM_switch_lp_conc_itm_7_1, or_tmp_21, NMP_RunFSM_switch_lp_conc_itm_7_2);
  assign NMP_PrepareReadReq_and_40_ssc = NMPRun_wen & (~ mux_13_nl) & and_dcpl_159
      & (~ NMP_RunFSM_switch_lp_conc_itm_7_3) & NMP_RunFSM_switch_lp_conc_itm_7_0;
  assign NMP_PrepareReadReq_and_68_enex5 = NMP_PrepareReadReq_and_40_ssc & reg_NMP_PrepareReadReq_asn_2_itm_6_enexo;
  assign NMP_PrepareWriteReq_and_83_enex5 = NMP_PrepareWriteReq_and_41_cse & reg_NMP_PrepareWriteReq_asn_1_itm_5_1_enexo_1;
  assign NMP_PrepareReadReq_and_69_enex5 = NMP_PrepareReadReq_and_44_cse & reg_NMP_PrepareReadReq_asn_2_itm_5_enexo;
  assign NMP_PrepareReadReq_and_70_enex5 = NMP_PrepareReadReq_and_44_cse & reg_NMP_PrepareReadReq_asn_2_itm_5_1_enexo_1;
  assign NMP_PrepareReadReq_and_71_enex5 = NMP_PrepareReadReq_and_44_cse & reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_2_enexo_1;
  assign and_880_nl = NMP_RunFSM_switch_lp_conc_itm_5_3 & NMP_RunFSM_switch_lp_conc_itm_5_1;
  assign mux_14_nl = MUX_s_1_2_2(and_880_nl, nor_58_cse, NMP_RunFSM_switch_lp_conc_itm_5_2);
  assign NMP_PrepareWriteReq_and_45_ssc = NMPRun_wen & mux_14_nl & and_dcpl_163 &
      (~ NMP_RunFSM_switch_lp_conc_itm_5_0);
  assign NMP_PrepareReadReq_and_72_enex5 = ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc
      & reg_NMP_PrepareReadReq_asn_2_itm_4_enexo;
  assign NMP_PrepareReadReq_and_48_ssc = NMPRun_wen & and_dcpl_166 & (~ NMP_RunFSM_switch_lp_conc_itm_4_1)
      & (~((~(NMP_RunFSM_switch_lp_conc_itm_4_2 ^ NMP_RunFSM_switch_lp_conc_itm_4_0))
      | NMP_RunFSM_switch_lp_conc_itm_4_3));
  assign out_adp_set_value_ac_float_1_and_12_ssc = NMPRun_wen & and_dcpl_554 & and_dcpl_557;
  assign out_adp_set_value_ac_float_1_and_13_ssc = NMPRun_wen & ((and_dcpl_564 &
      and_dcpl_567) | and_dcpl_509);
  assign out_adp_set_value_ac_float_1_and_14_ssc = NMPRun_wen & (state_2_sva ^ state_3_sva)
      & state_0_sva & (~(state_1_sva | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign rva_out_reg_data_and_5_ssc = NMPRun_wen & ((~ while_stage_0_3) | while_and_142_rgt)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign NMP_PrepareReadReq_and_73_enex5 = large_req_reg_write_data_data_and_64_cse
      & reg_NMP_PrepareReadReq_asn_1_itm_15_1_enexo;
  assign NMP_PrepareReadReq_and_74_enex5 = NMP_PrepareReadReq_and_17_cse & reg_NMP_PrepareReadReq_asn_1_itm_14_1_enexo;
  assign NMP_PrepareWriteReq_and_84_enex5 = NMP_PrepareWriteReq_and_24_cse & reg_NMP_PrepareWriteReq_asn_2_itm_11_enexo;
  assign NMP_PrepareWriteReq_and_85_enex5 = NMP_PrepareWriteReq_and_24_cse & reg_NMP_PrepareWriteReq_asn_2_itm_11_1_enexo;
  assign NMP_PrepareWriteReq_and_86_enex5 = NMP_PrepareWriteReq_and_24_cse & reg_NMP_PrepareWriteReq_asn_1_itm_11_2_enexo;
  assign out_adp_set_value_ac_float_1_and_4_ssc = NMPRun_wen & and_dcpl_101 & and_dcpl_105
      & NMP_RunFSM_switch_lp_conc_itm_12_0;
  assign out_adp_set_value_ac_float_and_4_ssc = NMPRun_wen & and_dcpl_101 & (~ NMP_RunFSM_switch_lp_conc_itm_12_3)
      & NMP_RunFSM_switch_lp_conc_itm_12_2 & NMP_RunFSM_switch_lp_conc_itm_12_0;
  assign NMP_PrepareReadReq_and_75_enex5 = NMP_PrepareReadReq_and_26_cse & reg_NMP_PrepareReadReq_asn_2_itm_11_enexo;
  assign NMP_PrepareReadReq_and_76_enex5 = NMP_PrepareReadReq_and_26_cse & reg_NMP_PrepareReadReq_asn_2_itm_11_1_enexo;
  assign NMP_PrepareWriteReq_and_27_ssc = NMPRun_wen & and_dcpl_124 & NMP_RunFSM_switch_lp_conc_itm_11_1
      & and_dcpl_130;
  assign NMP_PrepareWriteReq_and_87_enex5 = NMP_PrepareWriteReq_and_27_ssc & reg_NMP_PrepareWriteReq_asn_2_itm_10_enexo;
  assign NMP_PrepareWriteReq_and_88_enex5 = NMP_PrepareWriteReq_and_27_ssc & reg_NMP_PrepareWriteReq_asn_2_itm_10_1_enexo;
  assign NMP_PrepareReadReq_and_29_ssc = NMPRun_wen & and_dcpl_125 & (~(NMP_RunFSM_switch_lp_conc_itm_11_2
      | NMP_RunFSM_switch_lp_conc_itm_11_3)) & NMP_RunFSM_switch_lp_conc_itm_11_0;
  assign NMP_PrepareReadReq_and_77_enex5 = NMP_PrepareReadReq_and_29_ssc & reg_NMP_PrepareReadReq_asn_2_itm_10_1_enexo;
  assign out_adp_set_value_ac_float_1_and_9_ssc = NMPRun_wen & and_dcpl_305 & and_dcpl_519
      & NMP_RunFSM_switch_lp_conc_itm_6_3;
  assign out_adp_set_value_ac_float_1_and_10_ssc = NMPRun_wen & and_dcpl_354 & NMP_RunFSM_switch_lp_conc_itm_5_0
      & NMP_RunFSM_switch_lp_conc_itm_5_3 & (~ NMP_RunFSM_switch_lp_conc_itm_5_2);
  assign NMP_PrepareWriteReq_and_89_enex5 = NMP_PrepareWriteReq_and_35_cse & reg_NMP_PrepareWriteReq_asn_1_itm_8_2_enexo;
  assign NMP_PrepareReadReq_and_78_enex5 = NMP_PrepareReadReq_and_36_cse & reg_NMP_PrepareReadReq_asn_2_itm_8_enexo;
  assign NMP_PrepareReadReq_and_79_enex5 = NMP_PrepareReadReq_and_36_cse & reg_NMP_PrepareReadReq_asn_1_itm_8_2_enexo;
  assign NMP_PrepareWriteReq_and_90_enex5 = NMP_PrepareWriteReq_and_38_cse & reg_NMP_PrepareWriteReq_asn_1_itm_7_2_enexo;
  assign NMP_PrepareReadReq_and_80_enex5 = NMP_PrepareReadReq_and_39_cse & reg_NMP_PrepareReadReq_asn_2_itm_7_enexo;
  assign NMP_PrepareReadReq_and_81_enex5 = NMP_PrepareReadReq_and_39_cse & reg_NMP_PrepareReadReq_asn_1_itm_7_2_enexo;
  assign NMP_PrepareWriteReq_and_4_ssc = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[33:32]==2'b00)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareWriteReq_and_5_ssc = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[33:32]==2'b01)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareWriteReq_and_6_ssc = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[33:32]==2'b10)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareWriteReq_and_7_ssc = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[33:32]==2'b11)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareReadReq_and_7_ssc = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[33:32]==2'b01)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareWriteReq_and_91_enex5 = NMP_PrepareWriteReq_and_15_cse & reg_NMP_PrepareWriteReq_asn_2_itm_14_enexo;
  assign NMP_PrepareWriteReq_and_92_enex5 = NMP_PrepareWriteReq_and_15_cse & reg_NMP_PrepareWriteReq_asn_2_itm_14_1_enexo;
  assign NMP_PrepareWriteReq_and_93_enex5 = NMP_PrepareWriteReq_and_15_cse & reg_NMP_PrepareWriteReq_asn_1_itm_14_2_enexo;
  assign NMP_PrepareReadReq_and_82_enex5 = NMP_PrepareReadReq_and_17_cse & reg_NMP_PrepareReadReq_asn_2_itm_14_enexo;
  assign NMP_PrepareReadReq_and_83_enex5 = NMP_PrepareReadReq_and_17_cse & reg_NMP_PrepareReadReq_asn_2_itm_14_1_enexo;
  assign NMP_PrepareWriteReq_and_94_enex5 = NMP_PrepareWriteReq_and_18_cse & reg_NMP_PrepareWriteReq_asn_2_itm_13_enexo;
  assign NMP_PrepareWriteReq_and_95_enex5 = NMP_PrepareWriteReq_and_18_cse & reg_NMP_PrepareWriteReq_asn_2_itm_13_1_enexo;
  assign out_adp_set_value_ac_float_1_and_2_ssc = NMPRun_wen & and_dcpl_362 & and_dcpl_360
      & NMP_RunFSM_switch_lp_conc_itm_14_3;
  assign out_adp_set_value_ac_float_and_2_ssc = NMPRun_wen & and_dcpl_362 & NMP_RunFSM_switch_lp_conc_itm_14_0
      & NMP_RunFSM_switch_lp_conc_itm_14_2 & (~ NMP_RunFSM_switch_lp_conc_itm_14_3);
  assign NMP_PrepareReadReq_and_84_enex5 = NMP_PrepareReadReq_and_20_cse & reg_NMP_PrepareReadReq_asn_2_itm_13_1_enexo;
  assign NMP_PrepareWriteReq_and_96_enex5 = NMP_PrepareWriteReq_and_27_ssc & reg_NMP_PrepareWriteReq_asn_1_itm_10_2_enexo;
  assign NMP_PrepareReadReq_and_85_enex5 = NMP_PrepareReadReq_and_29_ssc & reg_NMP_PrepareReadReq_asn_2_itm_10_enexo;
  assign NMP_PrepareWriteReq_and_97_enex5 = NMP_PrepareWriteReq_and_21_cse & reg_NMP_PrepareWriteReq_asn_1_itm_12_2_enexo;
  assign NMP_PrepareReadReq_and_86_enex5 = NMP_PrepareReadReq_and_23_cse & reg_NMP_PrepareReadReq_asn_2_itm_12_enexo;
  assign NMP_PrepareWriteReq_and_98_enex5 = NMP_PrepareWriteReq_and_18_cse & reg_NMP_PrepareWriteReq_asn_1_itm_13_2_enexo;
  assign NMP_PrepareReadReq_and_87_enex5 = NMP_PrepareReadReq_and_20_cse & reg_NMP_PrepareReadReq_asn_2_itm_13_enexo;
  assign NMP_PrepareReadReq_and_88_enex5 = large_req_reg_write_data_data_and_64_cse
      & reg_NMP_PrepareReadReq_asn_2_itm_15_enexo;
  assign NMP_PrepareWriteReq_and_99_enex5 = NMP_PrepareWriteReq_and_12_cse & reg_NMP_PrepareWriteReq_asn_1_itm_15_2_enexo;
  assign out_float_round_32_if_m_1_and_15_tmp = NMPRun_wen & ((or_dcpl_110 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_31_tmp = NMPRun_wen & or_dcpl_110 & and_dcpl_177;
  assign out_float_round_32_1_if_m_1_and_31_tmp = NMPRun_wen & or_dcpl_222 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_15_tmp = NMPRun_wen & ((or_dcpl_222 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_14_tmp = NMPRun_wen & ((or_dcpl_103 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_30_tmp = NMPRun_wen & or_dcpl_103 & and_dcpl_177;
  assign out_float_round_32_1_if_m_1_and_14_tmp = NMPRun_wen & ((or_dcpl_215 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_30_tmp = NMPRun_wen & or_dcpl_215 & and_dcpl_195;
  assign out_float_round_32_if_m_1_and_29_tmp = NMPRun_wen & or_dcpl_96 & and_dcpl_177;
  assign out_float_round_32_if_m_1_and_13_tmp = NMPRun_wen & ((or_dcpl_96 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_29_tmp = NMPRun_wen & or_dcpl_208 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_13_tmp = NMPRun_wen & ((or_dcpl_208 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_12_tmp = NMPRun_wen & ((or_dcpl_89 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_28_tmp = NMPRun_wen & or_dcpl_89 & and_dcpl_177;
  assign out_float_round_32_1_if_m_1_and_12_tmp = NMPRun_wen & ((or_dcpl_201 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_28_tmp = NMPRun_wen & or_dcpl_201 & and_dcpl_195;
  assign out_float_round_32_if_m_1_and_27_tmp = NMPRun_wen & or_dcpl_82 & and_dcpl_177;
  assign out_float_round_32_if_m_1_and_11_tmp = NMPRun_wen & ((or_dcpl_82 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_27_tmp = NMPRun_wen & or_dcpl_194 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_11_tmp = NMPRun_wen & ((or_dcpl_194 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_26_tmp = NMPRun_wen & or_dcpl_75 & and_dcpl_177;
  assign out_float_round_32_if_m_1_and_10_tmp = NMPRun_wen & ((or_dcpl_75 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_10_tmp = NMPRun_wen & ((or_dcpl_187 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_26_tmp = NMPRun_wen & or_dcpl_187 & and_dcpl_195;
  assign out_float_round_32_if_m_1_and_25_tmp = NMPRun_wen & or_dcpl_68 & and_dcpl_177;
  assign out_float_round_32_if_m_1_and_9_tmp = NMPRun_wen & ((or_dcpl_68 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_25_tmp = NMPRun_wen & or_dcpl_180 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_9_tmp = NMPRun_wen & ((or_dcpl_180 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_24_tmp = NMPRun_wen & or_dcpl_61 & and_dcpl_177;
  assign out_float_round_32_if_m_1_and_8_tmp = NMPRun_wen & ((or_dcpl_61 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_8_tmp = NMPRun_wen & ((or_dcpl_173 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_24_tmp = NMPRun_wen & or_dcpl_173 & and_dcpl_195;
  assign out_float_round_32_if_m_1_and_7_tmp = NMPRun_wen & ((or_dcpl_54 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_23_tmp = NMPRun_wen & or_dcpl_54 & and_dcpl_177;
  assign out_float_round_32_1_if_m_1_and_23_tmp = NMPRun_wen & or_dcpl_166 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_7_tmp = NMPRun_wen & ((or_dcpl_166 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_22_tmp = NMPRun_wen & or_dcpl_47 & and_dcpl_177;
  assign out_float_round_32_if_m_1_and_6_tmp = NMPRun_wen & ((or_dcpl_47 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_22_tmp = NMPRun_wen & or_dcpl_159 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_6_tmp = NMPRun_wen & ((or_dcpl_159 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_21_tmp = NMPRun_wen & or_dcpl_40 & and_dcpl_177;
  assign out_float_round_32_if_m_1_and_5_tmp = NMPRun_wen & ((or_dcpl_40 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_21_tmp = NMPRun_wen & or_dcpl_152 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_5_tmp = NMPRun_wen & ((or_dcpl_152 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_20_tmp = NMPRun_wen & or_dcpl_33 & and_dcpl_177;
  assign out_float_round_32_if_m_1_and_4_tmp = NMPRun_wen & ((or_dcpl_33 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_4_tmp = NMPRun_wen & ((or_dcpl_145 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_20_tmp = NMPRun_wen & or_dcpl_145 & and_dcpl_195;
  assign out_float_round_32_if_m_1_and_19_tmp = NMPRun_wen & or_dcpl_26 & and_dcpl_177;
  assign out_float_round_32_if_m_1_and_3_tmp = NMPRun_wen & ((or_dcpl_26 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_19_tmp = NMPRun_wen & or_dcpl_138 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_3_tmp = NMPRun_wen & ((or_dcpl_138 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_2_tmp = NMPRun_wen & ((or_dcpl_19 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_18_tmp = NMPRun_wen & or_dcpl_19 & and_dcpl_177;
  assign out_float_round_32_1_if_m_1_and_18_tmp = NMPRun_wen & or_dcpl_131 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_2_tmp = NMPRun_wen & ((or_dcpl_131 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_1_tmp = NMPRun_wen & ((or_dcpl_12 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_17_tmp = NMPRun_wen & or_dcpl_12 & and_dcpl_177;
  assign out_float_round_32_1_if_m_1_and_1_tmp = NMPRun_wen & ((or_dcpl_124 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign out_float_round_32_1_if_m_1_and_17_tmp = NMPRun_wen & or_dcpl_124 & and_dcpl_195;
  assign out_float_round_32_if_m_1_and_tmp = NMPRun_wen & ((or_dcpl_5 & and_dcpl_10)
      | NMP_RunFSM_switch_lp_equal_tmp_4_15) & and_dcpl_5;
  assign out_float_round_32_if_m_1_and_16_tmp = NMPRun_wen & or_dcpl_5 & and_dcpl_177;
  assign out_float_round_32_1_if_m_1_and_16_tmp = NMPRun_wen & or_dcpl_117 & and_dcpl_195;
  assign out_float_round_32_1_if_m_1_and_tmp = NMPRun_wen & ((or_dcpl_117 & and_dcpl_47)
      | NMP_RunFSM_switch_lp_equal_tmp_8_15) & and_dcpl_5;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp = NMPRun_wen
      & (~ mux_tmp_7) & and_dcpl_283;
  assign NMP_ComputeSoftmaxMax_for_if_and_tmp = NMPRun_wen & and_dcpl_342;
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_tmp = NMPRun_wen
      & (~(((sum_exp_39_4_sva_st_2==36'b000000000000000000000000000000000000)) |
      or_dcpl_718 | NMP_RunFSM_switch_lp_conc_itm_10_2 | (~ NMP_RunFSM_switch_lp_conc_itm_10_3)
      | NMP_RunFSM_switch_lp_conc_itm_10_1 | NMP_RunFSM_switch_lp_conc_itm_10_0));
  assign and_1081_nl = ((~(state_0_sva | NMP_RunFSM_switch_lp_equal_tmp_10_1 | NMP_RunFSM_switch_lp_equal_tmp_11_1))
      | NMP_RunFSM_switch_lp_equal_tmp_1) & mux_cse;
  assign and_1080_nl = ((~((~ state_1_sva) | (~ state_0_sva) | NMP_RunFSM_switch_lp_equal_tmp_10_1
      | NMP_RunFSM_switch_lp_equal_tmp_11_1)) | NMP_RunFSM_switch_lp_equal_tmp_1)
      & mux_cse;
  assign mux_271_nl = MUX_s_1_2_2(and_1081_nl, and_1080_nl, state_3_sva);
  assign and_1079_nl = ((~((~ state_3_sva) | state_1_sva | state_0_sva | NMP_RunFSM_switch_lp_equal_tmp_10_1
      | NMP_RunFSM_switch_lp_equal_tmp_11_1)) | NMP_RunFSM_switch_lp_equal_tmp_1)
      & mux_cse;
  assign mux_272_nl = MUX_s_1_2_2(mux_271_nl, and_1079_nl, state_2_sva);
  assign nand_21_nl = ~(nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1
      & (~(NMP_RunFSM_switch_lp_equal_tmp_1 & mux_cse)));
  assign mux_273_nl = MUX_s_1_2_2(mux_272_nl, nand_21_nl, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign and_1082_tmp = mux_273_nl & NMPRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign or_976_nl = state_0_sva | (~ state_3_sva);
  assign mux_267_nl = MUX_s_1_2_2(or_534_cse, or_976_nl, state_2_sva);
  assign mux_266_nl = MUX_s_1_2_2(state_3_sva, (~ state_3_sva), state_0_sva);
  assign or_975_nl = state_2_sva | mux_266_nl;
  assign mux_268_nl = MUX_s_1_2_2(mux_267_nl, or_975_nl, state_1_sva);
  assign nor_294_nl = ~(NMP_RunFSM_switch_lp_equal_tmp_11_1 | NMP_RunFSM_switch_lp_equal_tmp_10_1
      | mux_268_nl);
  assign mux_269_nl = MUX_s_1_2_2(nor_294_nl, mux_cse, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign and_1063_tmp = (mux_269_nl | (NMP_RunFSM_switch_lp_equal_tmp_12_1 & (~ nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1)))
      & while_stage_0_3 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & NMPRun_wen;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo_ir_15_cse
          <= 1'b0;
      reg_NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo_ir_15_cse <= 1'b0;
      reg_NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo_ir_15_cse
          <= 1'b0;
      reg_NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo_ir_15_cse <= 1'b0;
      reg_done_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_large_rsp_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_large_req_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_4_39
          <= 1'b0;
      while_stage_0_3 <= 1'b0;
      while_stage_0_4 <= 1'b0;
      while_stage_0_5 <= 1'b0;
      while_stage_0_6 <= 1'b0;
      while_stage_0_7 <= 1'b0;
      while_stage_0_8 <= 1'b0;
      while_stage_0_9 <= 1'b0;
      while_stage_0_10 <= 1'b0;
      while_stage_0_11 <= 1'b0;
      while_stage_0_12 <= 1'b0;
      while_stage_0_13 <= 1'b0;
      while_stage_0_14 <= 1'b0;
      while_stage_0_15 <= 1'b0;
      while_stage_0_16 <= 1'b0;
      while_stage_0_17 <= 1'b0;
      while_stage_0_18 <= 1'b0;
      while_stage_0_19 <= 1'b0;
      while_stage_0_20 <= 1'b0;
      operator_3_false_operator_3_false_and_1_itm_2 <= 1'b0;
      operator_3_false_operator_3_false_and_1_itm_1 <= 1'b0;
      reg_NMP_PrepareReadReq_asn_1_itm_10_ftd <= 1'b0;
      reg_NMP_PrepareReadReq_asn_1_itm_10_ftd_1 <= 1'b0;
      NMP_PrepareReadReq_asn_1_itm_10_5_0 <= 6'b000000;
    end
    else if ( NMPRun_wen ) begin
      reg_NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_cgo_ir_15_cse
          <= and_582_rmff;
      reg_NMP_ComputeRMSNormalize_for_1_mul_cmp_cgo_ir_15_cse <= and_583_rmff;
      reg_NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_cgo_ir_15_cse
          <= and_584_rmff;
      reg_NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_cgo_ir_15_cse <= and_585_rmff;
      reg_done_Push_mioi_iswt0_cse <= and_587_rmff;
      reg_rva_out_Push_mioi_iswt0_cse <= and_588_rmff;
      reg_large_rsp_PopNB_mioi_iswt0_cse <= and_590_rmff;
      reg_start_PopNB_mioi_iswt0_cse <= and_591_rmff;
      reg_large_req_Push_mioi_iswt0_cse <= nor_206_rmff;
      reg_rva_in_PopNB_mioi_iswt0_cse <= fsm_output;
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_4_39
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_3_39;
      while_stage_0_3 <= reg_rva_in_PopNB_mioi_iswt0_cse;
      while_stage_0_4 <= while_stage_0_3;
      while_stage_0_5 <= while_stage_0_4;
      while_stage_0_6 <= while_stage_0_5;
      while_stage_0_7 <= while_stage_0_6;
      while_stage_0_8 <= while_stage_0_7;
      while_stage_0_9 <= while_stage_0_8;
      while_stage_0_10 <= while_stage_0_9;
      while_stage_0_11 <= while_stage_0_10;
      while_stage_0_12 <= while_stage_0_11;
      while_stage_0_13 <= while_stage_0_12;
      while_stage_0_14 <= while_stage_0_13;
      while_stage_0_15 <= while_stage_0_14;
      while_stage_0_16 <= while_stage_0_15;
      while_stage_0_17 <= while_stage_0_16;
      while_stage_0_18 <= while_stage_0_17;
      while_stage_0_19 <= while_stage_0_18;
      while_stage_0_20 <= while_stage_0_19;
      operator_3_false_operator_3_false_and_1_itm_2 <= operator_3_false_operator_3_false_and_1_itm_1;
      operator_3_false_operator_3_false_and_1_itm_1 <= (nmp_config_mode_sva_mx1==3'b001);
      reg_NMP_PrepareReadReq_asn_1_itm_10_ftd <= NMP_PrepareReadReq_asn_1_itm_9_rsp_0;
      reg_NMP_PrepareReadReq_asn_1_itm_10_ftd_1 <= NMP_PrepareReadReq_asn_1_itm_9_rsp_1_rsp_0;
      NMP_PrepareReadReq_asn_1_itm_10_5_0 <= MUX_v_6_2_2(NMP_PrepareReadReq_asn_1_itm_9_rsp_1_rsp_1,
          rtn_out, NMP_PrepareReadReq_or_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_1_mul_cmp_15_b_cse <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_13)
        & NMPRun_wen & or_928_cse & while_stage_0_15 ) begin
      reg_NMP_ComputeRMSNormalize_for_1_mul_cmp_15_b_cse <= rms_reciprocal_mux_rmff;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_b_cse <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_13)
        & NMPRun_wen & or_929_cse & while_stage_0_15 ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_b_cse <= sum_exp_reciprocal_mux_rmff;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      write_data_data_15_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_14_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_13_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_12_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_11_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_10_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_9_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_8_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_7_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_6_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_5_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_4_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_3_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_2_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_1_3_0_sva_dfm_1 <= 4'b0000;
      write_data_data_0_3_0_sva_dfm_1 <= 4'b0000;
    end
    else if ( and_936_cse ) begin
      write_data_data_15_3_0_sva_dfm_1 <= write_data_data_15_3_0_sva_dfm_1_mx0w0;
      write_data_data_14_3_0_sva_dfm_1 <= write_data_data_14_3_0_sva_dfm_1_mx0w0;
      write_data_data_13_3_0_sva_dfm_1 <= write_data_data_13_3_0_sva_dfm_1_mx0w0;
      write_data_data_12_3_0_sva_dfm_1 <= write_data_data_12_3_0_sva_dfm_1_mx0w0;
      write_data_data_11_3_0_sva_dfm_1 <= write_data_data_11_3_0_sva_dfm_1_mx0w0;
      write_data_data_10_3_0_sva_dfm_1 <= write_data_data_10_3_0_sva_dfm_1_mx0w0;
      write_data_data_9_3_0_sva_dfm_1 <= write_data_data_9_3_0_sva_dfm_1_mx0w0;
      write_data_data_8_3_0_sva_dfm_1 <= write_data_data_8_3_0_sva_dfm_1_mx0w0;
      write_data_data_7_3_0_sva_dfm_1 <= write_data_data_7_3_0_sva_dfm_1_mx0w0;
      write_data_data_6_3_0_sva_dfm_1 <= write_data_data_6_3_0_sva_dfm_1_mx0w0;
      write_data_data_5_3_0_sva_dfm_1 <= write_data_data_5_3_0_sva_dfm_1_mx0w0;
      write_data_data_4_3_0_sva_dfm_1 <= write_data_data_4_3_0_sva_dfm_1_mx0w0;
      write_data_data_3_3_0_sva_dfm_1 <= write_data_data_3_3_0_sva_dfm_1_mx0w0;
      write_data_data_2_3_0_sva_dfm_1 <= write_data_data_2_3_0_sva_dfm_1_mx0w0;
      write_data_data_1_3_0_sva_dfm_1 <= write_data_data_1_3_0_sva_dfm_1_mx0w0;
      write_data_data_0_3_0_sva_dfm_1 <= write_data_data_0_3_0_sva_dfm_1_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_16_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_16_nl,
          4'b1111, out_adp_set_value_ac_float_lor_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_16_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_16_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_15_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_17_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_15_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_17_nl,
          4'b1111, out_adp_set_value_ac_float_lor_15_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_15_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_17_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_15_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_17_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_15_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_14_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_18_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_14_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_18_nl,
          4'b1111, out_adp_set_value_ac_float_lor_14_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_14_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_18_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_14_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_18_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_14_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_13_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_19_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_13_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_19_nl,
          4'b1111, out_adp_set_value_ac_float_lor_13_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_13_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_19_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_13_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_19_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_13_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_12_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_20_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_12_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_20_nl,
          4'b1111, out_adp_set_value_ac_float_lor_12_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_12_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_20_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_12_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_20_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_12_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_11_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_21_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_11_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_21_nl,
          4'b1111, out_adp_set_value_ac_float_lor_11_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_11_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_21_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_11_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_21_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_11_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_10_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_22_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_10_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_22_nl,
          4'b1111, out_adp_set_value_ac_float_lor_10_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_10_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_22_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_10_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_22_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_10_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_9_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_23_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_9_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_23_nl,
          4'b1111, out_adp_set_value_ac_float_lor_9_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_9_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_23_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_9_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_23_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_9_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_8_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_24_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_8_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_24_nl,
          4'b1111, out_adp_set_value_ac_float_lor_8_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_8_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_24_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_8_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_24_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_8_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_7_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_25_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_7_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_25_nl,
          4'b1111, out_adp_set_value_ac_float_lor_7_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_7_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_25_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_7_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_25_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_7_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_6_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_26_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_6_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_26_nl,
          4'b1111, out_adp_set_value_ac_float_lor_6_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_6_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_26_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_6_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_26_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_6_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_5_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_27_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_5_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_27_nl,
          4'b1111, out_adp_set_value_ac_float_lor_5_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_5_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_27_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_5_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_27_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_5_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_4_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_28_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_4_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_28_nl,
          4'b1111, out_adp_set_value_ac_float_lor_4_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_4_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_28_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_4_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_28_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_4_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_3_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_29_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_3_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_29_nl,
          4'b1111, out_adp_set_value_ac_float_lor_3_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_3_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_29_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_3_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_29_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_3_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_2_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_30_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_2_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_30_nl,
          4'b1111, out_adp_set_value_ac_float_lor_2_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_2_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_30_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_2_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_30_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_2_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_1_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_31_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_for_out_adp_man_1_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_nor_31_nl,
          4'b1111, out_adp_set_value_ac_float_lor_1_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_1_lpi_1_dfm_1_1 <= 4'b0000;
    end
    else if ( NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_31_enex5 ) begin
      NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_1_lpi_1_dfm_1_1 <= ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_nor_31_nl,
          4'b1111, out_adp_set_value_ac_float_1_lor_1_lpi_1_dfm_1));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_equal_tmp_8_17 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_18
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_18 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_18 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_18 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_18 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_17 <= 1'b0;
      write_data_data_15_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_15_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_0_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_0_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_14_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_14_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_1_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_1_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_13_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_13_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_2_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_2_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_12_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_12_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_3_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_3_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_11_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_11_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_4_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_4_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_10_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_10_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_5_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_5_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_9_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_9_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_6_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_6_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_8_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_8_6_4_sva_dfm_1_0 <= 1'b0;
      write_data_data_7_6_4_sva_dfm_1_2_1 <= 2'b00;
      write_data_data_7_6_4_sva_dfm_1_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_cse ) begin
      NMP_RunFSM_switch_lp_equal_tmp_8_17 <= NMP_RunFSM_switch_lp_equal_tmp_8_16;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_18
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17;
      NMP_RunFSM_switch_lp_equal_tmp_4_17 <= NMP_RunFSM_switch_lp_equal_tmp_4_16;
      NMP_RunFSM_switch_lp_equal_tmp_18 <= NMP_RunFSM_switch_lp_equal_tmp_17_1;
      NMP_RunFSM_switch_lp_equal_tmp_1_17 <= NMP_RunFSM_switch_lp_equal_tmp_1_16;
      NMP_RunFSM_switch_lp_equal_tmp_2_17 <= NMP_RunFSM_switch_lp_equal_tmp_2_16;
      NMP_RunFSM_switch_lp_equal_tmp_3_17 <= NMP_RunFSM_switch_lp_equal_tmp_3_16;
      NMP_RunFSM_switch_lp_equal_tmp_5_17 <= NMP_RunFSM_switch_lp_equal_tmp_5_16;
      NMP_RunFSM_switch_lp_equal_tmp_6_17 <= NMP_RunFSM_switch_lp_equal_tmp_6_16;
      NMP_RunFSM_switch_lp_equal_tmp_7_17 <= NMP_RunFSM_switch_lp_equal_tmp_7_16;
      NMP_RunFSM_switch_lp_equal_tmp_9_17 <= NMP_RunFSM_switch_lp_equal_tmp_9_16;
      NMP_RunFSM_switch_lp_equal_tmp_10_18 <= NMP_RunFSM_switch_lp_equal_tmp_10_17;
      NMP_RunFSM_switch_lp_equal_tmp_11_18 <= NMP_RunFSM_switch_lp_equal_tmp_11_17;
      NMP_RunFSM_switch_lp_equal_tmp_12_18 <= NMP_RunFSM_switch_lp_equal_tmp_12_17;
      NMP_RunFSM_switch_lp_or_tmp_17 <= NMP_RunFSM_switch_lp_or_tmp_16;
      write_data_data_15_6_4_sva_dfm_1_2_1 <= write_data_data_15_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_15_6_4_sva_dfm_1_0 <= write_data_data_15_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_0_6_4_sva_dfm_1_2_1 <= write_data_data_0_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_0_6_4_sva_dfm_1_0 <= write_data_data_0_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_14_6_4_sva_dfm_1_2_1 <= write_data_data_14_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_14_6_4_sva_dfm_1_0 <= write_data_data_14_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_1_6_4_sva_dfm_1_2_1 <= write_data_data_1_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_1_6_4_sva_dfm_1_0 <= write_data_data_1_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_13_6_4_sva_dfm_1_2_1 <= write_data_data_13_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_13_6_4_sva_dfm_1_0 <= write_data_data_13_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_2_6_4_sva_dfm_1_2_1 <= write_data_data_2_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_2_6_4_sva_dfm_1_0 <= write_data_data_2_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_12_6_4_sva_dfm_1_2_1 <= write_data_data_12_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_12_6_4_sva_dfm_1_0 <= write_data_data_12_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_3_6_4_sva_dfm_1_2_1 <= write_data_data_3_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_3_6_4_sva_dfm_1_0 <= write_data_data_3_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_11_6_4_sva_dfm_1_2_1 <= write_data_data_11_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_11_6_4_sva_dfm_1_0 <= write_data_data_11_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_4_6_4_sva_dfm_1_2_1 <= write_data_data_4_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_4_6_4_sva_dfm_1_0 <= write_data_data_4_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_10_6_4_sva_dfm_1_2_1 <= write_data_data_10_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_10_6_4_sva_dfm_1_0 <= write_data_data_10_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_5_6_4_sva_dfm_1_2_1 <= write_data_data_5_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_5_6_4_sva_dfm_1_0 <= write_data_data_5_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_9_6_4_sva_dfm_1_2_1 <= write_data_data_9_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_9_6_4_sva_dfm_1_0 <= write_data_data_9_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_6_6_4_sva_dfm_1_2_1 <= write_data_data_6_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_6_6_4_sva_dfm_1_0 <= write_data_data_6_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_8_6_4_sva_dfm_1_2_1 <= write_data_data_8_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_8_6_4_sva_dfm_1_0 <= write_data_data_8_6_4_sva_dfm_1_0_mx0w0;
      write_data_data_7_6_4_sva_dfm_1_2_1 <= write_data_data_7_6_4_sva_dfm_1_2_1_mx0w0;
      write_data_data_7_6_4_sva_dfm_1_0 <= write_data_data_7_6_4_sva_dfm_1_0_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_req_reg_write_data_data_asn_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_1_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_1_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_46_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_46_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_45_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_3_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_4_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_4_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_43_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_43_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_42_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_6_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_7_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_7_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_40_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_40_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_39_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_9_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_10_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_10_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_37_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_37_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_36_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_12_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_13_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_13_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_34_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_34_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_33_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_15_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_16_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_16_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_31_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_31_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_30_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_18_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_19_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_19_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_28_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_28_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_27_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_21_itm_1 <= 1'b0;
      large_req_reg_write_data_data_asn_22_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_22_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_25_itm_1_2_1 <= 2'b00;
      large_req_reg_write_data_data_asn_25_itm_1_0 <= 1'b0;
      large_req_reg_write_data_data_asn_24_itm_1 <= 1'b0;
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_17 <= 2'b00;
      reg_NMP_PrepareReadReq_asn_1_itm_16_ftd <= 1'b0;
      reg_NMP_PrepareReadReq_asn_1_itm_16_ftd_1 <= 1'b0;
      reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_2_0 <= 3'b000;
    end
    else if ( large_req_reg_write_data_data_and_64_cse ) begin
      large_req_reg_write_data_data_asn_itm_1 <= large_req_reg_write_data_data_127_sva;
      large_req_reg_write_data_data_asn_1_itm_1_2_1 <= large_req_reg_write_data_data_126_124_sva_2_1;
      large_req_reg_write_data_data_asn_1_itm_1_0 <= large_req_reg_write_data_data_126_124_sva_0;
      large_req_reg_write_data_data_asn_46_itm_1_2_1 <= large_req_reg_write_data_data_6_4_sva_2_1;
      large_req_reg_write_data_data_asn_46_itm_1_0 <= large_req_reg_write_data_data_6_4_sva_0;
      large_req_reg_write_data_data_asn_45_itm_1 <= large_req_reg_write_data_data_7_sva;
      large_req_reg_write_data_data_asn_3_itm_1 <= large_req_reg_write_data_data_119_sva;
      large_req_reg_write_data_data_asn_4_itm_1_2_1 <= large_req_reg_write_data_data_118_116_sva_2_1;
      large_req_reg_write_data_data_asn_4_itm_1_0 <= large_req_reg_write_data_data_118_116_sva_0;
      large_req_reg_write_data_data_asn_43_itm_1_2_1 <= large_req_reg_write_data_data_14_12_sva_2_1;
      large_req_reg_write_data_data_asn_43_itm_1_0 <= large_req_reg_write_data_data_14_12_sva_0;
      large_req_reg_write_data_data_asn_42_itm_1 <= large_req_reg_write_data_data_15_sva;
      large_req_reg_write_data_data_asn_6_itm_1 <= large_req_reg_write_data_data_111_sva;
      large_req_reg_write_data_data_asn_7_itm_1_2_1 <= large_req_reg_write_data_data_110_108_sva_2_1;
      large_req_reg_write_data_data_asn_7_itm_1_0 <= large_req_reg_write_data_data_110_108_sva_0;
      large_req_reg_write_data_data_asn_40_itm_1_2_1 <= large_req_reg_write_data_data_22_20_sva_2_1;
      large_req_reg_write_data_data_asn_40_itm_1_0 <= large_req_reg_write_data_data_22_20_sva_0;
      large_req_reg_write_data_data_asn_39_itm_1 <= large_req_reg_write_data_data_23_sva;
      large_req_reg_write_data_data_asn_9_itm_1 <= large_req_reg_write_data_data_103_sva;
      large_req_reg_write_data_data_asn_10_itm_1_2_1 <= large_req_reg_write_data_data_102_100_sva_2_1;
      large_req_reg_write_data_data_asn_10_itm_1_0 <= large_req_reg_write_data_data_102_100_sva_0;
      large_req_reg_write_data_data_asn_37_itm_1_2_1 <= large_req_reg_write_data_data_30_28_sva_2_1;
      large_req_reg_write_data_data_asn_37_itm_1_0 <= large_req_reg_write_data_data_30_28_sva_0;
      large_req_reg_write_data_data_asn_36_itm_1 <= large_req_reg_write_data_data_31_sva;
      large_req_reg_write_data_data_asn_12_itm_1 <= large_req_reg_write_data_data_95_sva;
      large_req_reg_write_data_data_asn_13_itm_1_2_1 <= large_req_reg_write_data_data_94_92_sva_2_1;
      large_req_reg_write_data_data_asn_13_itm_1_0 <= large_req_reg_write_data_data_94_92_sva_0;
      large_req_reg_write_data_data_asn_34_itm_1_2_1 <= large_req_reg_write_data_data_38_36_sva_2_1;
      large_req_reg_write_data_data_asn_34_itm_1_0 <= large_req_reg_write_data_data_38_36_sva_0;
      large_req_reg_write_data_data_asn_33_itm_1 <= large_req_reg_write_data_data_39_sva;
      large_req_reg_write_data_data_asn_15_itm_1 <= large_req_reg_write_data_data_87_sva;
      large_req_reg_write_data_data_asn_16_itm_1_2_1 <= large_req_reg_write_data_data_86_84_sva_2_1;
      large_req_reg_write_data_data_asn_16_itm_1_0 <= large_req_reg_write_data_data_86_84_sva_0;
      large_req_reg_write_data_data_asn_31_itm_1_2_1 <= large_req_reg_write_data_data_46_44_sva_2_1;
      large_req_reg_write_data_data_asn_31_itm_1_0 <= large_req_reg_write_data_data_46_44_sva_0;
      large_req_reg_write_data_data_asn_30_itm_1 <= large_req_reg_write_data_data_47_sva;
      large_req_reg_write_data_data_asn_18_itm_1 <= large_req_reg_write_data_data_79_sva;
      large_req_reg_write_data_data_asn_19_itm_1_2_1 <= large_req_reg_write_data_data_78_76_sva_2_1;
      large_req_reg_write_data_data_asn_19_itm_1_0 <= large_req_reg_write_data_data_78_76_sva_0;
      large_req_reg_write_data_data_asn_28_itm_1_2_1 <= large_req_reg_write_data_data_54_52_sva_2_1;
      large_req_reg_write_data_data_asn_28_itm_1_0 <= large_req_reg_write_data_data_54_52_sva_0;
      large_req_reg_write_data_data_asn_27_itm_1 <= large_req_reg_write_data_data_55_sva;
      large_req_reg_write_data_data_asn_21_itm_1 <= large_req_reg_write_data_data_71_sva;
      large_req_reg_write_data_data_asn_22_itm_1_2_1 <= large_req_reg_write_data_data_70_68_sva_2_1;
      large_req_reg_write_data_data_asn_22_itm_1_0 <= large_req_reg_write_data_data_70_68_sva_0;
      large_req_reg_write_data_data_asn_25_itm_1_2_1 <= large_req_reg_write_data_data_62_60_sva_2_1;
      large_req_reg_write_data_data_asn_25_itm_1_0 <= large_req_reg_write_data_data_62_60_sva_0;
      large_req_reg_write_data_data_asn_24_itm_1 <= large_req_reg_write_data_data_63_sva;
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_17 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_16;
      reg_NMP_PrepareReadReq_asn_1_itm_16_ftd <= NMP_PrepareReadReq_asn_1_itm_15_7_6_rsp_0;
      reg_NMP_PrepareReadReq_asn_1_itm_16_ftd_1 <= NMP_PrepareReadReq_asn_1_itm_15_7_6_rsp_1;
      reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_2_0 <= reg_NMP_PrepareReadReq_asn_2_itm_15_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_req_reg_write_data_data_3_0_sva <= 4'b0000;
      large_req_reg_write_data_data_123_120_sva <= 4'b0000;
      large_req_reg_write_data_data_11_8_sva <= 4'b0000;
      large_req_reg_write_data_data_115_112_sva <= 4'b0000;
      large_req_reg_write_data_data_19_16_sva <= 4'b0000;
      large_req_reg_write_data_data_107_104_sva <= 4'b0000;
      large_req_reg_write_data_data_27_24_sva <= 4'b0000;
      large_req_reg_write_data_data_99_96_sva <= 4'b0000;
      large_req_reg_write_data_data_35_32_sva <= 4'b0000;
      large_req_reg_write_data_data_91_88_sva <= 4'b0000;
      large_req_reg_write_data_data_43_40_sva <= 4'b0000;
      large_req_reg_write_data_data_83_80_sva <= 4'b0000;
      large_req_reg_write_data_data_51_48_sva <= 4'b0000;
      large_req_reg_write_data_data_75_72_sva <= 4'b0000;
      large_req_reg_write_data_data_59_56_sva <= 4'b0000;
      large_req_reg_write_data_data_67_64_sva <= 4'b0000;
    end
    else if ( large_req_reg_write_data_data_and_cse ) begin
      large_req_reg_write_data_data_3_0_sva <= write_data_data_0_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_123_120_sva <= write_data_data_15_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_11_8_sva <= write_data_data_1_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_115_112_sva <= write_data_data_14_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_19_16_sva <= write_data_data_2_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_107_104_sva <= write_data_data_13_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_27_24_sva <= write_data_data_3_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_99_96_sva <= write_data_data_12_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_35_32_sva <= write_data_data_4_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_91_88_sva <= write_data_data_11_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_43_40_sva <= write_data_data_5_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_83_80_sva <= write_data_data_10_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_51_48_sva <= write_data_data_6_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_75_72_sva <= write_data_data_9_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_59_56_sva <= write_data_data_7_3_0_sva_dfm_1_mx1;
      large_req_reg_write_data_data_67_64_sva <= write_data_data_8_3_0_sva_dfm_1_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareReadReq_and_55_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_1 <= NMP_PrepareReadReq_asn_2_itm_15_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_3_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_tmp ) begin
      out_float_round_32_if_m_1_3_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_4_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_1_tmp ) begin
      out_float_round_32_if_m_1_4_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_5_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_2_tmp ) begin
      out_float_round_32_if_m_1_5_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_6_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_3_tmp ) begin
      out_float_round_32_if_m_1_6_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_7_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_4_tmp ) begin
      out_float_round_32_if_m_1_7_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_8_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_5_tmp ) begin
      out_float_round_32_if_m_1_8_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_9_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_6_tmp ) begin
      out_float_round_32_if_m_1_9_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_10_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_7_tmp ) begin
      out_float_round_32_if_m_1_10_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_11_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_8_tmp ) begin
      out_float_round_32_if_m_1_11_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_12_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_9_tmp ) begin
      out_float_round_32_if_m_1_12_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_13_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_10_tmp ) begin
      out_float_round_32_if_m_1_13_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_14_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_11_tmp ) begin
      out_float_round_32_if_m_1_14_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_15_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_12_tmp ) begin
      out_float_round_32_if_m_1_15_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_16_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_13_tmp ) begin
      out_float_round_32_if_m_1_16_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_17_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_14_tmp ) begin
      out_float_round_32_if_m_1_17_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_1_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_if_m_1_and_15_tmp ) begin
      out_float_round_32_if_m_1_1_sva_1_6 <= NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_16_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_15_itm_1
          <= 5'b00000;
      reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd <= 1'b0;
      reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1 <= 2'b00;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_14_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_14_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_13_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_13_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_12_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_11_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_10_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_9_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_9_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_8_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_7_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_7_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_6_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_5_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_4_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_4_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_3_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_3_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_2_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_2_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_1_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_itm_1
          <= 5'b00000;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse ) begin
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_16_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_sva_1 | (NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_15_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_30_nl);
      reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd <= out_adp_set_value_ac_float_asn_15_itm_15_rsp_0;
      reg_out_adp_set_value_ac_float_asn_15_itm_16_ftd_1 <= out_adp_set_value_ac_float_asn_15_itm_15_rsp_1;
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_15_sva_1 | (NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_14_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_29_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_14_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_14_sva_1 | (NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_13_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_28_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_13_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_13_sva_1 | (NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_12_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_27_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_12_sva_1 | (NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_11_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_26_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_11_sva_1 | (NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_10_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_25_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_10_sva_1 | (NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_9_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_24_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_9_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_9_sva_1 | (NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_8_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_23_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_8_sva_1 | (NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_7_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_22_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_7_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_7_sva_1 | (NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_6_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_21_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_6_sva_1 | (NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_5_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_20_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_5_sva_1 | (NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_4_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_19_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_4_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_4_sva_1 | (NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_3_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_18_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_3_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_3_sva_1 | (NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_2_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_17_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_2_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_2_sva_1 | (NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_1_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_16_nl);
      in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_for_out_float_m_4_1_sva_1 | (NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_3_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_tmp ) begin
      out_float_round_32_1_if_m_1_3_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_4_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_1_tmp ) begin
      out_float_round_32_1_if_m_1_4_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_5_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_2_tmp ) begin
      out_float_round_32_1_if_m_1_5_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_6_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_3_tmp ) begin
      out_float_round_32_1_if_m_1_6_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_7_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_4_tmp ) begin
      out_float_round_32_1_if_m_1_7_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_8_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_5_tmp ) begin
      out_float_round_32_1_if_m_1_8_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_9_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_6_tmp ) begin
      out_float_round_32_1_if_m_1_9_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_10_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_7_tmp ) begin
      out_float_round_32_1_if_m_1_10_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_11_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_8_tmp ) begin
      out_float_round_32_1_if_m_1_11_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_12_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_9_tmp ) begin
      out_float_round_32_1_if_m_1_12_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_13_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_10_tmp ) begin
      out_float_round_32_1_if_m_1_13_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_14_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_11_tmp ) begin
      out_float_round_32_1_if_m_1_14_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_15_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_12_tmp ) begin
      out_float_round_32_1_if_m_1_15_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_16_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_13_tmp ) begin
      out_float_round_32_1_if_m_1_16_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_17_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_14_tmp ) begin
      out_float_round_32_1_if_m_1_17_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_1_sva_1_6 <= 1'b0;
    end
    else if ( out_float_round_32_1_if_m_1_and_15_tmp ) begin
      out_float_round_32_1_if_m_1_1_sva_1_6 <= NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_16_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_15_itm_1
          <= 5'b00000;
      reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd <= 1'b0;
      reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1 <= 2'b00;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_15_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_14_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_13_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_13_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_12_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_12_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_11_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_11_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_10_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_9_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_9_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_8_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_7_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_7_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_6_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_5_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_5_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_4_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_3_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_2_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_1_itm_1
          <= 5'b00000;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1
          <= 1'b0;
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_itm_1
          <= 5'b00000;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse ) begin
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_16_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_15_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_30_nl);
      reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd <= out_adp_set_value_ac_float_1_asn_15_itm_15_rsp_0;
      reg_out_adp_set_value_ac_float_1_asn_15_itm_16_ftd_1 <= out_adp_set_value_ac_float_1_asn_15_itm_15_rsp_1;
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_15_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_15_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_14_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_29_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_14_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_13_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_28_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_13_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_13_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_12_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_27_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_12_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_12_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_11_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_26_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_11_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_11_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_10_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_25_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_10_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_9_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_24_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_9_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_9_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_8_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_23_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_8_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_7_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_22_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_7_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_7_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_6_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_21_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_6_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_5_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_20_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_5_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_5_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_4_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_19_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_4_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_3_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_18_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_3_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_2_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_17_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_2_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_1_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_16_nl);
      in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1
          <= ~((NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp[6])
          | NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_1_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000));
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_itm_1
          <= MUX_v_5_2_2(5'b00000, NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl,
          out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      write_data_data_15_7_sva_dfm_1 <= 1'b0;
      write_data_data_0_7_sva_dfm_1 <= 1'b0;
      write_data_data_14_7_sva_dfm_1 <= 1'b0;
      write_data_data_1_7_sva_dfm_1 <= 1'b0;
      write_data_data_13_7_sva_dfm_1 <= 1'b0;
      write_data_data_2_7_sva_dfm_1 <= 1'b0;
      write_data_data_12_7_sva_dfm_1 <= 1'b0;
      write_data_data_3_7_sva_dfm_1 <= 1'b0;
      write_data_data_11_7_sva_dfm_1 <= 1'b0;
      write_data_data_4_7_sva_dfm_1 <= 1'b0;
      write_data_data_10_7_sva_dfm_1 <= 1'b0;
      write_data_data_5_7_sva_dfm_1 <= 1'b0;
      write_data_data_9_7_sva_dfm_1 <= 1'b0;
      write_data_data_6_7_sva_dfm_1 <= 1'b0;
      write_data_data_8_7_sva_dfm_1 <= 1'b0;
      write_data_data_7_7_sva_dfm_1 <= 1'b0;
    end
    else if ( write_data_data_and_16_cse ) begin
      write_data_data_15_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_905_mx0w0;
      write_data_data_0_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_860_mx0w0;
      write_data_data_14_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_902_mx0w0;
      write_data_data_1_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_863_mx0w0;
      write_data_data_13_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_899_mx0w0;
      write_data_data_2_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_866_mx0w0;
      write_data_data_12_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_896_mx0w0;
      write_data_data_3_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_869_mx0w0;
      write_data_data_11_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_893_mx0w0;
      write_data_data_4_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_872_mx0w0;
      write_data_data_10_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_890_mx0w0;
      write_data_data_5_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_875_mx0w0;
      write_data_data_9_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_887_mx0w0;
      write_data_data_6_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_878_mx0w0;
      write_data_data_8_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_884_mx0w0;
      write_data_data_7_7_sva_dfm_1 <= NMP_RunFSM_switch_lp_mux1h_881_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_16_ftd <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_61_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_16_ftd <= NMP_PrepareWriteReq_asn_2_itm_15_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_16_ftd_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareWriteReq_and_62_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_16_ftd_1 <= NMP_PrepareWriteReq_asn_2_itm_15_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd <= 1'b0;
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_17 <= 2'b00;
      reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd_1_6 <= 1'b0;
    end
    else if ( NMP_PrepareWriteReq_and_12_cse ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd <= NMP_PrepareWriteReq_asn_1_itm_15_rsp_0;
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_17 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_16;
      reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd_1_6 <= reg_NMP_PrepareWriteReq_asn_1_itm_15_1_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_17_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_17_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_17_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_17_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_39_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_17_3 <= NMP_RunFSM_switch_lp_conc_itm_16_3;
      NMP_RunFSM_switch_lp_conc_itm_17_2 <= NMP_RunFSM_switch_lp_conc_itm_16_2;
      NMP_RunFSM_switch_lp_conc_itm_17_1 <= NMP_RunFSM_switch_lp_conc_itm_16_1;
      NMP_RunFSM_switch_lp_conc_itm_17_0 <= NMP_RunFSM_switch_lp_conc_itm_16_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_17 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_17_2 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_17_1_0 <= 2'b00;
      rva_out_reg_data_10_8_sva_dfm_3_17 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_17 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_6_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_17 <= rva_out_reg_data_0_sva_dfm_3_16;
      rva_out_reg_data_98_96_sva_dfm_3_17_2 <= reg_rva_out_reg_data_98_96_sva_dfm_3_16_ftd;
      rva_out_reg_data_98_96_sva_dfm_3_17_1_0 <= reg_rva_out_reg_data_98_96_sva_dfm_3_16_ftd_1;
      rva_out_reg_data_10_8_sva_dfm_3_17 <= rva_out_reg_data_10_8_sva_dfm_3_16;
      rva_out_reg_data_34_32_sva_dfm_3_17 <= rva_out_reg_data_34_32_sva_dfm_3_16;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_17 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_102_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_17 <= rva_out_reg_data_79_64_sva_dfm_3_16;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_17 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_103_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_17 <= rva_out_reg_data_55_48_sva_dfm_3_16;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_17 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ while_while_nor_itm_16) & while_stage_0_18 ) begin
      while_while_and_itm_17 <= while_while_and_itm_16;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_nor_itm_17 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_17_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_17 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_17 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_16 <= 1'b0;
    end
    else if ( while_and_144_cse ) begin
      while_while_nor_itm_17 <= while_while_nor_itm_16;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_17
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_16;
      NMP_RunFSM_switch_lp_equal_tmp_4_16 <= NMP_RunFSM_switch_lp_equal_tmp_4_15;
      NMP_RunFSM_switch_lp_equal_tmp_8_16 <= NMP_RunFSM_switch_lp_equal_tmp_8_15;
      NMP_RunFSM_switch_lp_equal_tmp_17_1 <= NMP_RunFSM_switch_lp_equal_tmp_16_1;
      NMP_RunFSM_switch_lp_equal_tmp_1_16 <= NMP_RunFSM_switch_lp_equal_tmp_1_15;
      NMP_RunFSM_switch_lp_equal_tmp_2_16 <= NMP_RunFSM_switch_lp_equal_tmp_2_15;
      NMP_RunFSM_switch_lp_equal_tmp_3_16 <= NMP_RunFSM_switch_lp_equal_tmp_3_15;
      NMP_RunFSM_switch_lp_equal_tmp_5_16 <= NMP_RunFSM_switch_lp_equal_tmp_5_15;
      NMP_RunFSM_switch_lp_equal_tmp_6_16 <= NMP_RunFSM_switch_lp_equal_tmp_6_15;
      NMP_RunFSM_switch_lp_equal_tmp_7_16 <= NMP_RunFSM_switch_lp_equal_tmp_7_15;
      NMP_RunFSM_switch_lp_equal_tmp_9_16 <= NMP_RunFSM_switch_lp_equal_tmp_9_15;
      NMP_RunFSM_switch_lp_equal_tmp_10_17 <= NMP_RunFSM_switch_lp_equal_tmp_10_16;
      NMP_RunFSM_switch_lp_equal_tmp_11_17 <= NMP_RunFSM_switch_lp_equal_tmp_11_16;
      NMP_RunFSM_switch_lp_equal_tmp_12_17 <= NMP_RunFSM_switch_lp_equal_tmp_12_16;
      NMP_RunFSM_switch_lp_or_tmp_16 <= NMP_RunFSM_switch_lp_or_tmp_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ComputeRMSNormalize_for_16_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_15_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_14_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_13_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_12_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_11_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_10_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_9_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_8_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_7_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_6_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_5_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_4_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_3_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_2_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeRMSNormalize_for_1_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      out_adp_set_value_ac_float_asn_15_itm_15_rsp_0 <= 1'b0;
      out_adp_set_value_ac_float_asn_15_itm_15_rsp_1 <= 2'b00;
    end
    else if ( out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_cse ) begin
      NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_out_2 & (~
          (NMP_ComputeRMSNormalize_for_1_mul_cmp_1_z[24]));
      NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_tmp;
      NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_out_2 & (~
          (NMP_ComputeRMSNormalize_for_1_mul_cmp_2_z[24]));
      NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_1_tmp;
      NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_out_2 & (~
          (NMP_ComputeRMSNormalize_for_1_mul_cmp_3_z[24]));
      NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_2_tmp;
      NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_out_2 & (~
          (NMP_ComputeRMSNormalize_for_1_mul_cmp_4_z[24]));
      NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_3_tmp;
      NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_out_2 & (~
          (NMP_ComputeRMSNormalize_for_1_mul_cmp_5_z[24]));
      NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_4_tmp;
      NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_out_2 & (~
          (NMP_ComputeRMSNormalize_for_1_mul_cmp_6_z[24]));
      NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_5_tmp;
      NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_out_2 & (~
          (NMP_ComputeRMSNormalize_for_1_mul_cmp_7_z[24]));
      NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_6_tmp;
      NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_out_2 & (~ (NMP_ComputeRMSNormalize_for_1_mul_cmp_8_z[24]));
      NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_7_tmp;
      NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_out_2 & (~ (NMP_ComputeRMSNormalize_for_1_mul_cmp_9_z[24]));
      NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_8_tmp;
      NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_out_2 & (~ (NMP_ComputeRMSNormalize_for_1_mul_cmp_10_z[24]));
      NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_9_tmp;
      NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_out_2 & (~ (NMP_ComputeRMSNormalize_for_1_mul_cmp_11_z[24]));
      NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_10_tmp;
      NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_out_2 & (~ (NMP_ComputeRMSNormalize_for_1_mul_cmp_12_z[24]));
      NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_11_tmp;
      NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_out_2 & (~ (NMP_ComputeRMSNormalize_for_1_mul_cmp_13_z[24]));
      NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_12_tmp;
      NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_out_2 & (~ (NMP_ComputeRMSNormalize_for_1_mul_cmp_14_z[24]));
      NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_13_tmp;
      NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_out_2 & (~ (NMP_ComputeRMSNormalize_for_1_mul_cmp_15_z[24]));
      NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_14_tmp;
      NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_out_2 & (~ (NMP_ComputeRMSNormalize_for_1_mul_cmp_z[24]));
      NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_15_tmp;
      NMP_ComputeRMSNormalize_for_16_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_1_z[55:24];
      NMP_ComputeRMSNormalize_for_15_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_2_z[55:24];
      NMP_ComputeRMSNormalize_for_14_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_3_z[55:24];
      NMP_ComputeRMSNormalize_for_13_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_4_z[55:24];
      NMP_ComputeRMSNormalize_for_12_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_5_z[55:24];
      NMP_ComputeRMSNormalize_for_11_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_6_z[55:24];
      NMP_ComputeRMSNormalize_for_10_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_7_z[55:24];
      NMP_ComputeRMSNormalize_for_9_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_8_z[55:24];
      NMP_ComputeRMSNormalize_for_8_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_9_z[55:24];
      NMP_ComputeRMSNormalize_for_7_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_10_z[55:24];
      NMP_ComputeRMSNormalize_for_6_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_11_z[55:24];
      NMP_ComputeRMSNormalize_for_5_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_12_z[55:24];
      NMP_ComputeRMSNormalize_for_4_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_13_z[55:24];
      NMP_ComputeRMSNormalize_for_3_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_14_z[55:24];
      NMP_ComputeRMSNormalize_for_2_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_15_z[55:24];
      NMP_ComputeRMSNormalize_for_1_slc_55_24_ncse_sva_1 <= NMP_ComputeRMSNormalize_for_1_mul_cmp_z[55:24];
      out_adp_set_value_ac_float_asn_15_itm_15_rsp_0 <= out_adp_set_value_ac_float_asn_15_itm_14_2;
      out_adp_set_value_ac_float_asn_15_itm_15_rsp_1 <= out_adp_set_value_ac_float_asn_15_itm_14_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= 1'b0;
      NMP_ComputeSoftmaxNormalize_for_16_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_15_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_14_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_13_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_12_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_11_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_10_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_9_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_8_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_7_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_6_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_5_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_4_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_3_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_2_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      NMP_ComputeSoftmaxNormalize_for_1_slc_55_24_ncse_sva_1 <= 32'b00000000000000000000000000000000;
      out_adp_set_value_ac_float_1_asn_15_itm_15_rsp_0 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_15_rsp_1 <= 2'b00;
    end
    else if ( out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_cse ) begin
      NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_1_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_2_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_3_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_4_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_5_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_6_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_7_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_8_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_9_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_10_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_11_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_12_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_13_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_14_tmp;
      NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1
          <= NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_out_2 &
          (~ (NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_z[24]));
      NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1
          <= out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_15_tmp;
      NMP_ComputeSoftmaxNormalize_for_16_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_15_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_14_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_13_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_12_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_11_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_10_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_9_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_8_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_7_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_6_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_5_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_4_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_3_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_2_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_z[55:24];
      NMP_ComputeSoftmaxNormalize_for_1_slc_55_24_ncse_sva_1 <= NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_z[55:24];
      out_adp_set_value_ac_float_1_asn_15_itm_15_rsp_0 <= out_adp_set_value_ac_float_1_asn_15_itm_14_2;
      out_adp_set_value_ac_float_1_asn_15_itm_15_rsp_1 <= out_adp_set_value_ac_float_1_asn_15_itm_14_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_16_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_16_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_16_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_16_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_43_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_16_3 <= NMP_RunFSM_switch_lp_conc_itm_15_3;
      NMP_RunFSM_switch_lp_conc_itm_16_2 <= NMP_RunFSM_switch_lp_conc_itm_15_2;
      NMP_RunFSM_switch_lp_conc_itm_16_1 <= NMP_RunFSM_switch_lp_conc_itm_15_1;
      NMP_RunFSM_switch_lp_conc_itm_16_0 <= NMP_RunFSM_switch_lp_conc_itm_15_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_16
          <= 1'b0;
      while_while_nor_itm_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_16 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_16 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_16_1 <= 1'b0;
    end
    else if ( while_if_and_2_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_16
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_15;
      while_while_nor_itm_16 <= while_while_nor_itm_15;
      NMP_RunFSM_switch_lp_equal_tmp_9_15 <= NMP_RunFSM_switch_lp_equal_tmp_9_14;
      NMP_RunFSM_switch_lp_equal_tmp_1_15 <= NMP_RunFSM_switch_lp_equal_tmp_1_14;
      NMP_RunFSM_switch_lp_equal_tmp_2_15 <= NMP_RunFSM_switch_lp_equal_tmp_2_14;
      NMP_RunFSM_switch_lp_equal_tmp_3_15 <= NMP_RunFSM_switch_lp_equal_tmp_3_14;
      NMP_RunFSM_switch_lp_equal_tmp_4_15 <= NMP_RunFSM_switch_lp_equal_tmp_4_14;
      NMP_RunFSM_switch_lp_equal_tmp_5_15 <= NMP_RunFSM_switch_lp_equal_tmp_5_14;
      NMP_RunFSM_switch_lp_equal_tmp_6_15 <= NMP_RunFSM_switch_lp_equal_tmp_6_14;
      NMP_RunFSM_switch_lp_equal_tmp_7_15 <= NMP_RunFSM_switch_lp_equal_tmp_7_14;
      NMP_RunFSM_switch_lp_equal_tmp_8_15 <= NMP_RunFSM_switch_lp_equal_tmp_8_14;
      NMP_RunFSM_switch_lp_equal_tmp_10_16 <= NMP_RunFSM_switch_lp_equal_tmp_10_15;
      NMP_RunFSM_switch_lp_equal_tmp_11_16 <= NMP_RunFSM_switch_lp_equal_tmp_11_15;
      NMP_RunFSM_switch_lp_equal_tmp_12_16 <= NMP_RunFSM_switch_lp_equal_tmp_12_15;
      NMP_RunFSM_switch_lp_or_tmp_15 <= NMP_RunFSM_switch_lp_or_tmp_14;
      NMP_RunFSM_switch_lp_equal_tmp_16_1 <= NMP_RunFSM_switch_lp_equal_tmp_15_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_15_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_15_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_15_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_15_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_47_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_15_3 <= NMP_RunFSM_switch_lp_conc_itm_14_3;
      NMP_RunFSM_switch_lp_conc_itm_15_2 <= NMP_RunFSM_switch_lp_conc_itm_14_2;
      NMP_RunFSM_switch_lp_conc_itm_15_1 <= NMP_RunFSM_switch_lp_conc_itm_14_1;
      NMP_RunFSM_switch_lp_conc_itm_15_0 <= NMP_RunFSM_switch_lp_conc_itm_14_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_15
          <= 1'b0;
      while_while_nor_itm_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_15 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_15 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_15_1 <= 1'b0;
    end
    else if ( while_if_and_3_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_15
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_14;
      while_while_nor_itm_15 <= while_while_nor_itm_14;
      NMP_RunFSM_switch_lp_equal_tmp_1_14 <= NMP_RunFSM_switch_lp_equal_tmp_1_13;
      NMP_RunFSM_switch_lp_equal_tmp_2_14 <= NMP_RunFSM_switch_lp_equal_tmp_2_13;
      NMP_RunFSM_switch_lp_equal_tmp_3_14 <= NMP_RunFSM_switch_lp_equal_tmp_3_13;
      NMP_RunFSM_switch_lp_equal_tmp_4_14 <= NMP_RunFSM_switch_lp_equal_tmp_4_13;
      NMP_RunFSM_switch_lp_equal_tmp_5_14 <= NMP_RunFSM_switch_lp_equal_tmp_5_13;
      NMP_RunFSM_switch_lp_equal_tmp_6_14 <= NMP_RunFSM_switch_lp_equal_tmp_6_13;
      NMP_RunFSM_switch_lp_equal_tmp_7_14 <= NMP_RunFSM_switch_lp_equal_tmp_7_13;
      NMP_RunFSM_switch_lp_equal_tmp_8_14 <= NMP_RunFSM_switch_lp_equal_tmp_8_13;
      NMP_RunFSM_switch_lp_equal_tmp_9_14 <= NMP_RunFSM_switch_lp_equal_tmp_9_13;
      NMP_RunFSM_switch_lp_equal_tmp_10_15 <= NMP_RunFSM_switch_lp_equal_tmp_10_14;
      NMP_RunFSM_switch_lp_equal_tmp_11_15 <= NMP_RunFSM_switch_lp_equal_tmp_11_14;
      NMP_RunFSM_switch_lp_equal_tmp_12_15 <= NMP_RunFSM_switch_lp_equal_tmp_12_14;
      NMP_RunFSM_switch_lp_or_tmp_14 <= NMP_RunFSM_switch_lp_or_tmp_13;
      NMP_RunFSM_switch_lp_equal_tmp_15_1 <= NMP_RunFSM_switch_lp_equal_tmp_14_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_14_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_14_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_14_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_14_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_51_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_14_3 <= NMP_RunFSM_switch_lp_conc_itm_13_3;
      NMP_RunFSM_switch_lp_conc_itm_14_2 <= NMP_RunFSM_switch_lp_conc_itm_13_2;
      NMP_RunFSM_switch_lp_conc_itm_14_1 <= NMP_RunFSM_switch_lp_conc_itm_13_1;
      NMP_RunFSM_switch_lp_conc_itm_14_0 <= NMP_RunFSM_switch_lp_conc_itm_13_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_14
          <= 1'b0;
      while_while_nor_itm_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_14 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_14 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_14_1 <= 1'b0;
    end
    else if ( while_if_and_4_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_14
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_13;
      while_while_nor_itm_14 <= while_while_nor_itm_13;
      NMP_RunFSM_switch_lp_equal_tmp_1_13 <= NMP_RunFSM_switch_lp_equal_tmp_1_12;
      NMP_RunFSM_switch_lp_equal_tmp_2_13 <= NMP_RunFSM_switch_lp_equal_tmp_2_12;
      NMP_RunFSM_switch_lp_equal_tmp_3_13 <= NMP_RunFSM_switch_lp_equal_tmp_3_12;
      NMP_RunFSM_switch_lp_equal_tmp_4_13 <= NMP_RunFSM_switch_lp_equal_tmp_4_12;
      NMP_RunFSM_switch_lp_equal_tmp_5_13 <= NMP_RunFSM_switch_lp_equal_tmp_5_12;
      NMP_RunFSM_switch_lp_equal_tmp_6_13 <= NMP_RunFSM_switch_lp_equal_tmp_6_12;
      NMP_RunFSM_switch_lp_equal_tmp_7_13 <= NMP_RunFSM_switch_lp_equal_tmp_7_12;
      NMP_RunFSM_switch_lp_equal_tmp_8_13 <= NMP_RunFSM_switch_lp_equal_tmp_8_12;
      NMP_RunFSM_switch_lp_equal_tmp_9_13 <= NMP_RunFSM_switch_lp_equal_tmp_9_12;
      NMP_RunFSM_switch_lp_equal_tmp_10_14 <= NMP_RunFSM_switch_lp_equal_tmp_10_13;
      NMP_RunFSM_switch_lp_equal_tmp_11_14 <= NMP_RunFSM_switch_lp_equal_tmp_11_13;
      NMP_RunFSM_switch_lp_equal_tmp_12_14 <= NMP_RunFSM_switch_lp_equal_tmp_12_13;
      NMP_RunFSM_switch_lp_or_tmp_13 <= NMP_RunFSM_switch_lp_or_tmp_12;
      NMP_RunFSM_switch_lp_equal_tmp_14_1 <= NMP_RunFSM_switch_lp_equal_tmp_13_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1_9_0
          <= 10'b0000000000;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5
        ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1_9_0
          <= MUX_v_10_2_2((ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_mx0w0[9:0]),
          ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_9_0,
          and_dcpl_634);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_3
          <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_3_enex5
        ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_3
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_3 <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_1_enex5
        ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_3 <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_equal_tmp_3_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_13_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_12 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_13
          <= 1'b0;
      while_while_nor_itm_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_13 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_13 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_12 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_55_cse ) begin
      NMP_RunFSM_switch_lp_equal_tmp_3_12 <= NMP_RunFSM_switch_lp_equal_tmp_3_11;
      NMP_RunFSM_switch_lp_equal_tmp_13_1 <= NMP_RunFSM_switch_lp_equal_tmp_12;
      NMP_RunFSM_switch_lp_equal_tmp_7_12 <= NMP_RunFSM_switch_lp_equal_tmp_7_11;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_13
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_12;
      while_while_nor_itm_13 <= while_while_nor_itm_12;
      NMP_RunFSM_switch_lp_equal_tmp_1_12 <= NMP_RunFSM_switch_lp_equal_tmp_1_11;
      NMP_RunFSM_switch_lp_equal_tmp_2_12 <= NMP_RunFSM_switch_lp_equal_tmp_2_11;
      NMP_RunFSM_switch_lp_equal_tmp_4_12 <= NMP_RunFSM_switch_lp_equal_tmp_4_11;
      NMP_RunFSM_switch_lp_equal_tmp_5_12 <= NMP_RunFSM_switch_lp_equal_tmp_5_11;
      NMP_RunFSM_switch_lp_equal_tmp_6_12 <= NMP_RunFSM_switch_lp_equal_tmp_6_11;
      NMP_RunFSM_switch_lp_equal_tmp_8_12 <= NMP_RunFSM_switch_lp_equal_tmp_8_11;
      NMP_RunFSM_switch_lp_equal_tmp_9_12 <= NMP_RunFSM_switch_lp_equal_tmp_9_11;
      NMP_RunFSM_switch_lp_equal_tmp_10_13 <= NMP_RunFSM_switch_lp_equal_tmp_10_12;
      NMP_RunFSM_switch_lp_equal_tmp_11_13 <= NMP_RunFSM_switch_lp_equal_tmp_11_12;
      NMP_RunFSM_switch_lp_equal_tmp_12_13 <= NMP_RunFSM_switch_lp_equal_tmp_12_12;
      NMP_RunFSM_switch_lp_or_tmp_12 <= NMP_RunFSM_switch_lp_or_tmp_11;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_4
          <= 1'b0;
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_5
          <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_56_cse ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_4
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_3;
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_5
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_13_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_13_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_13_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_13_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_60_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_13_3 <= NMP_RunFSM_switch_lp_conc_itm_12_3;
      NMP_RunFSM_switch_lp_conc_itm_13_2 <= NMP_RunFSM_switch_lp_conc_itm_12_2;
      NMP_RunFSM_switch_lp_conc_itm_13_1 <= NMP_RunFSM_switch_lp_conc_itm_12_1;
      NMP_RunFSM_switch_lp_conc_itm_13_0 <= NMP_RunFSM_switch_lp_conc_itm_12_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_3
          <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_3
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_145_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_10 <= NMP_ComputeRMSNormalize_for_asn_60_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_146_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_10 <= NMP_ComputeRMSNormalize_for_asn_58_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_147_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_10 <= NMP_ComputeRMSNormalize_for_asn_56_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_148_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_10 <= NMP_ComputeRMSNormalize_for_asn_54_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_149_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_10 <= NMP_ComputeRMSNormalize_for_asn_52_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_150_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_10 <= NMP_ComputeRMSNormalize_for_asn_50_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_151_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_10 <= NMP_ComputeRMSNormalize_for_asn_48_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_152_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_10 <= NMP_ComputeRMSNormalize_for_asn_46_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_153_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_10 <= NMP_ComputeRMSNormalize_for_asn_44_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_154_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_10 <= NMP_ComputeRMSNormalize_for_asn_42_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_155_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_10 <= NMP_ComputeRMSNormalize_for_asn_40_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_156_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_10 <= NMP_ComputeRMSNormalize_for_asn_38_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_157_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_10 <= NMP_ComputeRMSNormalize_for_asn_36_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_11 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_158_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_11 <= NMP_ComputeRMSNormalize_for_asn_34_itm_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_11 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_159_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_11 <= NMP_ComputeRMSNormalize_for_asn_32_itm_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_11 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_160_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_11 <= NMP_ComputeRMSNormalize_for_asn_itm_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      sum_exp_39_4_sva_st_4 <= 36'b000000000000000000000000000000000000;
    end
    else if ( sum_exp_and_enex5 ) begin
      sum_exp_39_4_sva_st_4 <= sum_exp_39_4_sva_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_45_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_80_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_45_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_45_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_43_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_81_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_43_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_43_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_41_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_82_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_41_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_41_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_39_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_83_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_39_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_39_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_37_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_84_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_37_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_37_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_35_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_85_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_35_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_35_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_33_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_86_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_33_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_33_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_31_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_87_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_31_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_31_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_29_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_88_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_29_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_29_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_27_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_89_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_27_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_27_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_25_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_90_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_25_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_25_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_23_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_91_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_23_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_23_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_21_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_92_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_21_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_21_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_19_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_93_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_19_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_19_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_17_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_94_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_17_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_17_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_itm_4 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_95_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_itm_4 <= NMP_ComputeSoftmaxNormalize_for_asn_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_12_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_12_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_12_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_12_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_64_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_12_3 <= NMP_RunFSM_switch_lp_conc_itm_11_3;
      NMP_RunFSM_switch_lp_conc_itm_12_2 <= NMP_RunFSM_switch_lp_conc_itm_11_2;
      NMP_RunFSM_switch_lp_conc_itm_12_1 <= NMP_RunFSM_switch_lp_conc_itm_11_1;
      NMP_RunFSM_switch_lp_conc_itm_12_0 <= NMP_RunFSM_switch_lp_conc_itm_11_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_12
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12 <= 1'b0;
      while_while_nor_itm_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_12 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_12 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_11 <= 1'b0;
    end
    else if ( while_if_and_6_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_12
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11;
      NMP_RunFSM_switch_lp_equal_tmp_3_11 <= NMP_RunFSM_switch_lp_equal_tmp_3_10;
      NMP_RunFSM_switch_lp_equal_tmp_7_11 <= NMP_RunFSM_switch_lp_equal_tmp_7_10;
      NMP_RunFSM_switch_lp_equal_tmp_12 <= NMP_RunFSM_switch_lp_equal_tmp_11;
      while_while_nor_itm_12 <= while_while_nor_itm_11;
      NMP_RunFSM_switch_lp_equal_tmp_1_11 <= NMP_RunFSM_switch_lp_equal_tmp_1_10;
      NMP_RunFSM_switch_lp_equal_tmp_2_11 <= NMP_RunFSM_switch_lp_equal_tmp_2_10;
      NMP_RunFSM_switch_lp_equal_tmp_4_11 <= NMP_RunFSM_switch_lp_equal_tmp_4_10;
      NMP_RunFSM_switch_lp_equal_tmp_5_11 <= NMP_RunFSM_switch_lp_equal_tmp_5_10;
      NMP_RunFSM_switch_lp_equal_tmp_6_11 <= NMP_RunFSM_switch_lp_equal_tmp_6_10;
      NMP_RunFSM_switch_lp_equal_tmp_8_11 <= NMP_RunFSM_switch_lp_equal_tmp_8_10;
      NMP_RunFSM_switch_lp_equal_tmp_9_11 <= NMP_RunFSM_switch_lp_equal_tmp_9_10;
      NMP_RunFSM_switch_lp_equal_tmp_10_12 <= NMP_RunFSM_switch_lp_equal_tmp_10_11;
      NMP_RunFSM_switch_lp_equal_tmp_11_12 <= NMP_RunFSM_switch_lp_equal_tmp_11_11;
      NMP_RunFSM_switch_lp_equal_tmp_12_12 <= NMP_RunFSM_switch_lp_equal_tmp_12_11;
      NMP_RunFSM_switch_lp_or_tmp_11 <= NMP_RunFSM_switch_lp_or_tmp_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_2
          <= 40'b0000000000000000000000000000000000000000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_1_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_2
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      sum_exp_39_4_sva_st_3 <= 36'b000000000000000000000000000000000000;
    end
    else if ( sum_exp_and_1_enex5 ) begin
      sum_exp_39_4_sva_st_3 <= sum_exp_39_4_sva_st_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_11_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_11_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_11_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_11_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_68_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_11_3 <= NMP_RunFSM_switch_lp_conc_itm_10_3;
      NMP_RunFSM_switch_lp_conc_itm_11_2 <= NMP_RunFSM_switch_lp_conc_itm_10_2;
      NMP_RunFSM_switch_lp_conc_itm_11_1 <= NMP_RunFSM_switch_lp_conc_itm_10_1;
      NMP_RunFSM_switch_lp_conc_itm_11_0 <= NMP_RunFSM_switch_lp_conc_itm_10_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11 <= 1'b0;
      while_while_nor_itm_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_11 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_11 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_10 <= 1'b0;
    end
    else if ( while_if_and_7_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10;
      NMP_RunFSM_switch_lp_equal_tmp_3_10 <= NMP_RunFSM_switch_lp_equal_tmp_3_9;
      NMP_RunFSM_switch_lp_equal_tmp_7_10 <= NMP_RunFSM_switch_lp_equal_tmp_7_9;
      NMP_RunFSM_switch_lp_equal_tmp_11 <= NMP_RunFSM_switch_lp_equal_tmp_10;
      while_while_nor_itm_11 <= while_while_nor_itm_10;
      NMP_RunFSM_switch_lp_equal_tmp_1_10 <= NMP_RunFSM_switch_lp_equal_tmp_1_9;
      NMP_RunFSM_switch_lp_equal_tmp_2_10 <= NMP_RunFSM_switch_lp_equal_tmp_2_9;
      NMP_RunFSM_switch_lp_equal_tmp_4_10 <= NMP_RunFSM_switch_lp_equal_tmp_4_9;
      NMP_RunFSM_switch_lp_equal_tmp_5_10 <= NMP_RunFSM_switch_lp_equal_tmp_5_9;
      NMP_RunFSM_switch_lp_equal_tmp_6_10 <= NMP_RunFSM_switch_lp_equal_tmp_6_9;
      NMP_RunFSM_switch_lp_equal_tmp_8_10 <= NMP_RunFSM_switch_lp_equal_tmp_8_9;
      NMP_RunFSM_switch_lp_equal_tmp_9_10 <= NMP_RunFSM_switch_lp_equal_tmp_9_9;
      NMP_RunFSM_switch_lp_equal_tmp_10_11 <= NMP_RunFSM_switch_lp_equal_tmp_10_10;
      NMP_RunFSM_switch_lp_equal_tmp_11_11 <= NMP_RunFSM_switch_lp_equal_tmp_11_10;
      NMP_RunFSM_switch_lp_equal_tmp_12_11 <= NMP_RunFSM_switch_lp_equal_tmp_12_10;
      NMP_RunFSM_switch_lp_or_tmp_10 <= NMP_RunFSM_switch_lp_or_tmp_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_1
          <= 40'b0000000000000000000000000000000000000000;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_39
          <= 1'b0;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_38_0
          <= 39'b000000000000000000000000000000000000000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_2_cse
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_1
          <= operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_39
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_mx0_39;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_38_0
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_mx0_38_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      sum_exp_39_4_sva_st_2 <= 36'b000000000000000000000000000000000000;
    end
    else if ( sum_exp_and_2_enex5 ) begin
      sum_exp_39_4_sva_st_2 <= sum_exp_39_4_sva_st_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_10_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_10_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_10_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_10_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_72_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_10_3 <= NMP_RunFSM_switch_lp_conc_itm_9_3;
      NMP_RunFSM_switch_lp_conc_itm_10_2 <= NMP_RunFSM_switch_lp_conc_itm_9_2;
      NMP_RunFSM_switch_lp_conc_itm_10_1 <= NMP_RunFSM_switch_lp_conc_itm_9_1;
      NMP_RunFSM_switch_lp_conc_itm_10_0 <= NMP_RunFSM_switch_lp_conc_itm_9_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10 <= 1'b0;
      while_while_nor_itm_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_10 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_10 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_9 <= 1'b0;
    end
    else if ( while_if_and_8_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
      NMP_RunFSM_switch_lp_equal_tmp_3_9 <= NMP_RunFSM_switch_lp_equal_tmp_3_8;
      NMP_RunFSM_switch_lp_equal_tmp_7_9 <= NMP_RunFSM_switch_lp_equal_tmp_7_8;
      NMP_RunFSM_switch_lp_equal_tmp_10 <= NMP_RunFSM_switch_lp_equal_tmp_9;
      while_while_nor_itm_10 <= while_while_nor_itm_9;
      NMP_RunFSM_switch_lp_equal_tmp_1_9 <= NMP_RunFSM_switch_lp_equal_tmp_1_8;
      NMP_RunFSM_switch_lp_equal_tmp_2_9 <= NMP_RunFSM_switch_lp_equal_tmp_2_8;
      NMP_RunFSM_switch_lp_equal_tmp_4_9 <= NMP_RunFSM_switch_lp_equal_tmp_4_8;
      NMP_RunFSM_switch_lp_equal_tmp_5_9 <= NMP_RunFSM_switch_lp_equal_tmp_5_8;
      NMP_RunFSM_switch_lp_equal_tmp_6_9 <= NMP_RunFSM_switch_lp_equal_tmp_6_8;
      NMP_RunFSM_switch_lp_equal_tmp_8_9 <= NMP_RunFSM_switch_lp_equal_tmp_8_8;
      NMP_RunFSM_switch_lp_equal_tmp_9_9 <= NMP_RunFSM_switch_lp_equal_tmp_9_8;
      NMP_RunFSM_switch_lp_equal_tmp_10_10 <= NMP_RunFSM_switch_lp_equal_tmp_10_9;
      NMP_RunFSM_switch_lp_equal_tmp_11_10 <= NMP_RunFSM_switch_lp_equal_tmp_11_9;
      NMP_RunFSM_switch_lp_equal_tmp_12_10 <= NMP_RunFSM_switch_lp_equal_tmp_12_9;
      NMP_RunFSM_switch_lp_or_tmp_9 <= NMP_RunFSM_switch_lp_or_tmp_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_itm_1
          <= 1'b0;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_2_cse
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_itm_1
          <= (ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_itm_35_11_1[0])
          & (ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4[0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_6_1_itm_1
          <= 6'b000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_12_enex5
        ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_6_1_itm_1
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4[6:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_9_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_9_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_9_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_9_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_76_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_9_3 <= NMP_RunFSM_switch_lp_conc_itm_8_3;
      NMP_RunFSM_switch_lp_conc_itm_9_2 <= NMP_RunFSM_switch_lp_conc_itm_8_2;
      NMP_RunFSM_switch_lp_conc_itm_9_1 <= NMP_RunFSM_switch_lp_conc_itm_8_1;
      NMP_RunFSM_switch_lp_conc_itm_9_0 <= NMP_RunFSM_switch_lp_conc_itm_8_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9 <= 1'b0;
      while_while_nor_itm_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_9 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_9 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_8 <= 1'b0;
    end
    else if ( while_if_and_9_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
      NMP_RunFSM_switch_lp_equal_tmp_3_8 <= NMP_RunFSM_switch_lp_equal_tmp_3_7;
      NMP_RunFSM_switch_lp_equal_tmp_7_8 <= NMP_RunFSM_switch_lp_equal_tmp_7_7;
      NMP_RunFSM_switch_lp_equal_tmp_9 <= NMP_RunFSM_switch_lp_equal_tmp_8;
      while_while_nor_itm_9 <= while_while_nor_itm_8;
      NMP_RunFSM_switch_lp_equal_tmp_1_8 <= NMP_RunFSM_switch_lp_equal_tmp_1_7;
      NMP_RunFSM_switch_lp_equal_tmp_2_8 <= NMP_RunFSM_switch_lp_equal_tmp_2_7;
      NMP_RunFSM_switch_lp_equal_tmp_4_8 <= NMP_RunFSM_switch_lp_equal_tmp_4_7;
      NMP_RunFSM_switch_lp_equal_tmp_5_8 <= NMP_RunFSM_switch_lp_equal_tmp_5_7;
      NMP_RunFSM_switch_lp_equal_tmp_6_8 <= NMP_RunFSM_switch_lp_equal_tmp_6_7;
      NMP_RunFSM_switch_lp_equal_tmp_8_8 <= NMP_RunFSM_switch_lp_equal_tmp_8_7;
      NMP_RunFSM_switch_lp_equal_tmp_9_8 <= NMP_RunFSM_switch_lp_equal_tmp_9_7;
      NMP_RunFSM_switch_lp_equal_tmp_10_9 <= NMP_RunFSM_switch_lp_equal_tmp_10_8;
      NMP_RunFSM_switch_lp_equal_tmp_11_9 <= NMP_RunFSM_switch_lp_equal_tmp_11_8;
      NMP_RunFSM_switch_lp_equal_tmp_12_9 <= NMP_RunFSM_switch_lp_equal_tmp_12_8;
      NMP_RunFSM_switch_lp_or_tmp_8 <= NMP_RunFSM_switch_lp_or_tmp_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_8_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_8_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_8_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_8_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_80_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_8_3 <= NMP_RunFSM_switch_lp_conc_itm_7_3;
      NMP_RunFSM_switch_lp_conc_itm_8_2 <= NMP_RunFSM_switch_lp_conc_itm_7_2;
      NMP_RunFSM_switch_lp_conc_itm_8_1 <= NMP_RunFSM_switch_lp_conc_itm_7_1;
      NMP_RunFSM_switch_lp_conc_itm_8_0 <= NMP_RunFSM_switch_lp_conc_itm_7_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_7 <= 1'b0;
      while_while_nor_itm_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_8 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_8 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_7 <= 1'b0;
    end
    else if ( while_if_and_10_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
      NMP_RunFSM_switch_lp_equal_tmp_6_7 <= NMP_RunFSM_switch_lp_equal_tmp_6_6;
      NMP_RunFSM_switch_lp_equal_tmp_8 <= NMP_RunFSM_switch_lp_equal_tmp_7;
      NMP_RunFSM_switch_lp_equal_tmp_3_7 <= NMP_RunFSM_switch_lp_equal_tmp_3_6;
      NMP_RunFSM_switch_lp_equal_tmp_7_7 <= NMP_RunFSM_switch_lp_equal_tmp_7_6;
      while_while_nor_itm_8 <= while_while_nor_itm_7;
      NMP_RunFSM_switch_lp_equal_tmp_1_7 <= NMP_RunFSM_switch_lp_equal_tmp_1_6;
      NMP_RunFSM_switch_lp_equal_tmp_2_7 <= NMP_RunFSM_switch_lp_equal_tmp_2_6;
      NMP_RunFSM_switch_lp_equal_tmp_4_7 <= NMP_RunFSM_switch_lp_equal_tmp_4_6;
      NMP_RunFSM_switch_lp_equal_tmp_5_7 <= NMP_RunFSM_switch_lp_equal_tmp_5_6;
      NMP_RunFSM_switch_lp_equal_tmp_8_7 <= NMP_RunFSM_switch_lp_equal_tmp_8_6;
      NMP_RunFSM_switch_lp_equal_tmp_9_7 <= NMP_RunFSM_switch_lp_equal_tmp_9_6;
      NMP_RunFSM_switch_lp_equal_tmp_10_8 <= NMP_RunFSM_switch_lp_equal_tmp_10_7;
      NMP_RunFSM_switch_lp_equal_tmp_11_8 <= NMP_RunFSM_switch_lp_equal_tmp_11_7;
      NMP_RunFSM_switch_lp_equal_tmp_12_8 <= NMP_RunFSM_switch_lp_equal_tmp_12_7;
      NMP_RunFSM_switch_lp_or_tmp_7 <= NMP_RunFSM_switch_lp_or_tmp_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_7_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_7_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_7_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_7_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_84_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_7_3 <= NMP_RunFSM_switch_lp_conc_itm_6_3;
      NMP_RunFSM_switch_lp_conc_itm_7_2 <= NMP_RunFSM_switch_lp_conc_itm_6_2;
      NMP_RunFSM_switch_lp_conc_itm_7_1 <= NMP_RunFSM_switch_lp_conc_itm_6_1;
      NMP_RunFSM_switch_lp_conc_itm_7_0 <= NMP_RunFSM_switch_lp_conc_itm_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_6 <= 1'b0;
      while_while_nor_itm_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_7 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_7 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_6 <= 1'b0;
    end
    else if ( while_if_and_11_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
      NMP_RunFSM_switch_lp_equal_tmp_6_6 <= NMP_RunFSM_switch_lp_equal_tmp_6_5;
      NMP_RunFSM_switch_lp_equal_tmp_7 <= NMP_RunFSM_switch_lp_equal_tmp_6;
      NMP_RunFSM_switch_lp_equal_tmp_3_6 <= NMP_RunFSM_switch_lp_equal_tmp_3_5;
      NMP_RunFSM_switch_lp_equal_tmp_7_6 <= NMP_RunFSM_switch_lp_equal_tmp_7_5;
      while_while_nor_itm_7 <= while_while_nor_itm_6;
      NMP_RunFSM_switch_lp_equal_tmp_1_6 <= NMP_RunFSM_switch_lp_equal_tmp_1_5;
      NMP_RunFSM_switch_lp_equal_tmp_2_6 <= NMP_RunFSM_switch_lp_equal_tmp_2_5;
      NMP_RunFSM_switch_lp_equal_tmp_4_6 <= NMP_RunFSM_switch_lp_equal_tmp_4_5;
      NMP_RunFSM_switch_lp_equal_tmp_5_6 <= NMP_RunFSM_switch_lp_equal_tmp_5_5;
      NMP_RunFSM_switch_lp_equal_tmp_8_6 <= NMP_RunFSM_switch_lp_equal_tmp_8_5;
      NMP_RunFSM_switch_lp_equal_tmp_9_6 <= NMP_RunFSM_switch_lp_equal_tmp_9_5;
      NMP_RunFSM_switch_lp_equal_tmp_10_7 <= NMP_RunFSM_switch_lp_equal_tmp_10_6;
      NMP_RunFSM_switch_lp_equal_tmp_11_7 <= NMP_RunFSM_switch_lp_equal_tmp_11_6;
      NMP_RunFSM_switch_lp_equal_tmp_12_7 <= NMP_RunFSM_switch_lp_equal_tmp_12_6;
      NMP_RunFSM_switch_lp_or_tmp_6 <= NMP_RunFSM_switch_lp_or_tmp_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_6_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_6_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_6_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_6_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_88_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_6_3 <= NMP_RunFSM_switch_lp_conc_itm_5_3;
      NMP_RunFSM_switch_lp_conc_itm_6_2 <= NMP_RunFSM_switch_lp_conc_itm_5_2;
      NMP_RunFSM_switch_lp_conc_itm_6_1 <= NMP_RunFSM_switch_lp_conc_itm_5_1;
      NMP_RunFSM_switch_lp_conc_itm_6_0 <= NMP_RunFSM_switch_lp_conc_itm_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_5 <= 1'b0;
      while_while_nor_itm_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_6 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_6 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_5 <= 1'b0;
    end
    else if ( while_if_and_12_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
      NMP_RunFSM_switch_lp_equal_tmp_6_5 <= NMP_RunFSM_switch_lp_equal_tmp_6_4;
      NMP_RunFSM_switch_lp_equal_tmp_6 <= NMP_RunFSM_switch_lp_equal_tmp_5;
      NMP_RunFSM_switch_lp_equal_tmp_3_5 <= NMP_RunFSM_switch_lp_equal_tmp_3_4;
      NMP_RunFSM_switch_lp_equal_tmp_7_5 <= NMP_RunFSM_switch_lp_equal_tmp_7_4;
      while_while_nor_itm_6 <= while_while_nor_itm_5;
      NMP_RunFSM_switch_lp_equal_tmp_1_5 <= NMP_RunFSM_switch_lp_equal_tmp_1_4;
      NMP_RunFSM_switch_lp_equal_tmp_2_5 <= NMP_RunFSM_switch_lp_equal_tmp_2_4;
      NMP_RunFSM_switch_lp_equal_tmp_4_5 <= NMP_RunFSM_switch_lp_equal_tmp_4_4;
      NMP_RunFSM_switch_lp_equal_tmp_5_5 <= NMP_RunFSM_switch_lp_equal_tmp_5_4;
      NMP_RunFSM_switch_lp_equal_tmp_8_5 <= NMP_RunFSM_switch_lp_equal_tmp_8_4;
      NMP_RunFSM_switch_lp_equal_tmp_9_5 <= NMP_RunFSM_switch_lp_equal_tmp_9_4;
      NMP_RunFSM_switch_lp_equal_tmp_10_6 <= NMP_RunFSM_switch_lp_equal_tmp_10_5;
      NMP_RunFSM_switch_lp_equal_tmp_11_6 <= NMP_RunFSM_switch_lp_equal_tmp_11_5;
      NMP_RunFSM_switch_lp_equal_tmp_12_6 <= NMP_RunFSM_switch_lp_equal_tmp_12_5;
      NMP_RunFSM_switch_lp_or_tmp_5 <= NMP_RunFSM_switch_lp_or_tmp_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_16_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_50_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_16_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_16_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_15_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_51_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_15_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_15_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_14_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_52_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_14_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_14_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_13_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_53_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_13_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_13_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_12_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_54_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_12_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_12_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_11_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_55_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_11_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_11_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_10_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_56_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_10_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_10_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_9_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_57_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_9_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_9_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_8_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_58_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_8_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_8_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_7_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_59_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_7_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_7_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_6_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_60_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_6_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_6_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_5_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_61_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_5_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_5_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_4_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_62_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_4_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_4_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_3_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_63_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_3_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_3_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_2_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_64_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_2_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_2_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_1_acc_1_itm_1 <= 28'b0000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_65_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_1_acc_1_itm_1 <= nl_NMP_ComputeSoftmaxExp_for_1_acc_1_itm_1[27:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_5_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_5_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_5_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_5_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_92_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_5_3 <= NMP_RunFSM_switch_lp_conc_itm_4_3;
      NMP_RunFSM_switch_lp_conc_itm_5_2 <= NMP_RunFSM_switch_lp_conc_itm_4_2;
      NMP_RunFSM_switch_lp_conc_itm_5_1 <= NMP_RunFSM_switch_lp_conc_itm_4_1;
      NMP_RunFSM_switch_lp_conc_itm_5_0 <= NMP_RunFSM_switch_lp_conc_itm_4_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_4 <= 1'b0;
      while_while_nor_itm_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_5 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_5 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_4 <= 1'b0;
    end
    else if ( while_if_and_13_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
      NMP_RunFSM_switch_lp_equal_tmp_5_4 <= NMP_RunFSM_switch_lp_equal_tmp_5_3;
      NMP_RunFSM_switch_lp_equal_tmp_5 <= NMP_RunFSM_switch_lp_equal_tmp_4;
      NMP_RunFSM_switch_lp_equal_tmp_6_4 <= NMP_RunFSM_switch_lp_equal_tmp_6_3;
      NMP_RunFSM_switch_lp_equal_tmp_3_4 <= NMP_RunFSM_switch_lp_equal_tmp_3_3;
      NMP_RunFSM_switch_lp_equal_tmp_7_4 <= NMP_RunFSM_switch_lp_equal_tmp_7_3;
      while_while_nor_itm_5 <= while_while_nor_itm_4;
      NMP_RunFSM_switch_lp_equal_tmp_1_4 <= NMP_RunFSM_switch_lp_equal_tmp_1_3;
      NMP_RunFSM_switch_lp_equal_tmp_2_4 <= NMP_RunFSM_switch_lp_equal_tmp_2_3;
      NMP_RunFSM_switch_lp_equal_tmp_4_4 <= NMP_RunFSM_switch_lp_equal_tmp_4_3;
      NMP_RunFSM_switch_lp_equal_tmp_8_4 <= NMP_RunFSM_switch_lp_equal_tmp_8_3;
      NMP_RunFSM_switch_lp_equal_tmp_9_4 <= NMP_RunFSM_switch_lp_equal_tmp_9_3;
      NMP_RunFSM_switch_lp_equal_tmp_10_5 <= NMP_RunFSM_switch_lp_equal_tmp_10_4;
      NMP_RunFSM_switch_lp_equal_tmp_11_5 <= NMP_RunFSM_switch_lp_equal_tmp_11_4;
      NMP_RunFSM_switch_lp_equal_tmp_12_5 <= NMP_RunFSM_switch_lp_equal_tmp_12_4;
      NMP_RunFSM_switch_lp_or_tmp_4 <= NMP_RunFSM_switch_lp_or_tmp_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_4_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_4_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_4_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_4_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_96_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_4_3 <= NMP_RunFSM_switch_lp_conc_itm_3_3;
      NMP_RunFSM_switch_lp_conc_itm_4_2 <= NMP_RunFSM_switch_lp_conc_itm_3_2;
      NMP_RunFSM_switch_lp_conc_itm_4_1 <= NMP_RunFSM_switch_lp_conc_itm_3_1;
      NMP_RunFSM_switch_lp_conc_itm_4_0 <= NMP_RunFSM_switch_lp_conc_itm_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_3 <= 1'b0;
      while_while_nor_itm_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_4 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_4 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_3 <= 1'b0;
    end
    else if ( while_if_and_14_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_3;
      NMP_RunFSM_switch_lp_equal_tmp_5_3 <= NMP_RunFSM_switch_lp_equal_tmp_5_2;
      NMP_RunFSM_switch_lp_equal_tmp_4 <= NMP_RunFSM_switch_lp_equal_tmp_3;
      NMP_RunFSM_switch_lp_equal_tmp_2_3 <= NMP_RunFSM_switch_lp_equal_tmp_2_2;
      NMP_RunFSM_switch_lp_equal_tmp_6_3 <= NMP_RunFSM_switch_lp_equal_tmp_6_2;
      NMP_RunFSM_switch_lp_equal_tmp_3_3 <= NMP_RunFSM_switch_lp_equal_tmp_3_2;
      NMP_RunFSM_switch_lp_equal_tmp_7_3 <= NMP_RunFSM_switch_lp_equal_tmp_7_2;
      while_while_nor_itm_4 <= while_while_nor_itm_3;
      NMP_RunFSM_switch_lp_equal_tmp_1_3 <= NMP_RunFSM_switch_lp_equal_tmp_1_2;
      NMP_RunFSM_switch_lp_equal_tmp_4_3 <= NMP_RunFSM_switch_lp_equal_tmp_4_2;
      NMP_RunFSM_switch_lp_equal_tmp_8_3 <= NMP_RunFSM_switch_lp_equal_tmp_8_2;
      NMP_RunFSM_switch_lp_equal_tmp_9_3 <= NMP_RunFSM_switch_lp_equal_tmp_9_2;
      NMP_RunFSM_switch_lp_equal_tmp_10_4 <= NMP_RunFSM_switch_lp_equal_tmp_10_3;
      NMP_RunFSM_switch_lp_equal_tmp_11_4 <= NMP_RunFSM_switch_lp_equal_tmp_11_3;
      NMP_RunFSM_switch_lp_equal_tmp_12_4 <= NMP_RunFSM_switch_lp_equal_tmp_12_3;
      NMP_RunFSM_switch_lp_or_tmp_3 <= NMP_RunFSM_switch_lp_or_tmp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_3_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_3_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_3_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_3_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_100_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_3_3 <= NMP_RunFSM_switch_lp_conc_itm_2_3;
      NMP_RunFSM_switch_lp_conc_itm_3_2 <= NMP_RunFSM_switch_lp_conc_itm_2_2;
      NMP_RunFSM_switch_lp_conc_itm_3_1 <= NMP_RunFSM_switch_lp_conc_itm_2_1;
      NMP_RunFSM_switch_lp_conc_itm_3_0 <= NMP_RunFSM_switch_lp_conc_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_3
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_2 <= 1'b0;
      while_while_nor_itm_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_3 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_3 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_2 <= 1'b0;
    end
    else if ( while_if_and_15_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_3
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
      NMP_RunFSM_switch_lp_equal_tmp_5_2 <= NMP_RunFSM_switch_lp_equal_tmp_5_1;
      NMP_RunFSM_switch_lp_equal_tmp_3 <= NMP_RunFSM_switch_lp_equal_tmp_2;
      NMP_RunFSM_switch_lp_equal_tmp_2_2 <= NMP_RunFSM_switch_lp_equal_tmp_2_1;
      NMP_RunFSM_switch_lp_equal_tmp_6_2 <= NMP_RunFSM_switch_lp_equal_tmp_6_1;
      NMP_RunFSM_switch_lp_equal_tmp_3_2 <= NMP_RunFSM_switch_lp_equal_tmp_3_1;
      NMP_RunFSM_switch_lp_equal_tmp_7_2 <= NMP_RunFSM_switch_lp_equal_tmp_7_1;
      while_while_nor_itm_3 <= while_while_nor_itm_2;
      NMP_RunFSM_switch_lp_equal_tmp_1_2 <= NMP_RunFSM_switch_lp_equal_tmp_1_1;
      NMP_RunFSM_switch_lp_equal_tmp_4_2 <= NMP_RunFSM_switch_lp_equal_tmp_4_1;
      NMP_RunFSM_switch_lp_equal_tmp_8_2 <= NMP_RunFSM_switch_lp_equal_tmp_8_1;
      NMP_RunFSM_switch_lp_equal_tmp_9_2 <= NMP_RunFSM_switch_lp_equal_tmp_9_1;
      NMP_RunFSM_switch_lp_equal_tmp_10_3 <= NMP_RunFSM_switch_lp_equal_tmp_10_2;
      NMP_RunFSM_switch_lp_equal_tmp_11_3 <= NMP_RunFSM_switch_lp_equal_tmp_11_2;
      NMP_RunFSM_switch_lp_equal_tmp_12_3 <= NMP_RunFSM_switch_lp_equal_tmp_12_2;
      NMP_RunFSM_switch_lp_or_tmp_2 <= NMP_RunFSM_switch_lp_or_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_fixed_15_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_14_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_13_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_12_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_11_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_10_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_9_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_8_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_7_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_6_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_5_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_4_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_3_26_0_sva <= 27'b000000000000000000000000000;
    end
    else if ( and_983_cse ) begin
      input_fixed_15_26_0_sva <= input_fixed_mux_7_cse;
      input_fixed_14_26_0_sva <= input_fixed_mux_5_cse;
      input_fixed_13_26_0_sva <= input_fixed_mux_3_cse;
      input_fixed_12_26_0_sva <= input_fixed_mux_1_cse;
      input_fixed_11_26_0_sva <= input_fixed_mux_25_cse;
      input_fixed_10_26_0_sva <= input_fixed_mux_23_cse;
      input_fixed_9_26_0_sva <= input_fixed_mux_21_cse;
      input_fixed_8_26_0_sva <= input_fixed_mux_19_cse;
      input_fixed_7_26_0_sva <= input_fixed_mux_17_cse;
      input_fixed_6_26_0_sva <= input_fixed_mux_15_cse;
      input_fixed_5_26_0_sva <= input_fixed_mux_13_cse;
      input_fixed_4_26_0_sva <= input_fixed_mux_11_cse;
      input_fixed_3_26_0_sva <= input_fixed_mux_9_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_conc_itm_2_3 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_2_2 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_2_1 <= 1'b0;
      NMP_RunFSM_switch_lp_conc_itm_2_0 <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_104_cse ) begin
      NMP_RunFSM_switch_lp_conc_itm_2_3 <= state_3_sva;
      NMP_RunFSM_switch_lp_conc_itm_2_2 <= state_2_sva;
      NMP_RunFSM_switch_lp_conc_itm_2_1 <= state_1_sva;
      NMP_RunFSM_switch_lp_conc_itm_2_0 <= state_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_fixed_15_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_14_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_13_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_12_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_11_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_10_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_9_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_8_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_7_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_6_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_5_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_4_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
      input_fixed_3_26_0_sva_dfm_2_1 <= 27'b000000000000000000000000000;
    end
    else if ( and_1011_cse ) begin
      input_fixed_15_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_51_nl,
          input_fixed_mux_7_cse, or_1057_cse);
      input_fixed_14_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_50_nl,
          input_fixed_mux_5_cse, or_1057_cse);
      input_fixed_13_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_49_nl,
          input_fixed_mux_3_cse, or_1057_cse);
      input_fixed_12_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_48_nl,
          input_fixed_mux_1_cse, or_1057_cse);
      input_fixed_11_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_47_nl,
          input_fixed_mux_25_cse, or_1057_cse);
      input_fixed_10_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_46_nl,
          input_fixed_mux_23_cse, or_1057_cse);
      input_fixed_9_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_45_nl,
          input_fixed_mux_21_cse, or_1057_cse);
      input_fixed_8_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_44_nl,
          input_fixed_mux_19_cse, or_1057_cse);
      input_fixed_7_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_43_nl,
          input_fixed_mux_17_cse, or_1057_cse);
      input_fixed_6_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_42_nl,
          input_fixed_mux_15_cse, or_1057_cse);
      input_fixed_5_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_41_nl,
          input_fixed_mux_13_cse, or_1057_cse);
      input_fixed_4_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_40_nl,
          input_fixed_mux_11_cse, or_1057_cse);
      input_fixed_3_26_0_sva_dfm_2_1 <= MUX_v_27_2_2(NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_39_nl,
          input_fixed_mux_9_cse, or_1057_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_5_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_2_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_6_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_3_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_7_1 <= 1'b0;
      while_while_nor_itm_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_4_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_8_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_9_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_2 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_2 <= 1'b0;
      NMP_RunFSM_switch_lp_or_tmp_1_1 <= 1'b0;
    end
    else if ( input_fixed_and_16_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
      NMP_RunFSM_switch_lp_equal_tmp_5_1 <= NMP_RunFSM_switch_lp_equal_tmp_17;
      NMP_RunFSM_switch_lp_equal_tmp_2 <= NMP_RunFSM_switch_lp_equal_tmp_1;
      NMP_RunFSM_switch_lp_equal_tmp_2_1 <= NMP_RunFSM_switch_lp_equal_tmp_18_1;
      NMP_RunFSM_switch_lp_equal_tmp_6_1 <= NMP_RunFSM_switch_lp_equal_tmp_19;
      NMP_RunFSM_switch_lp_equal_tmp_3_1 <= NMP_RunFSM_switch_lp_equal_tmp_20;
      NMP_RunFSM_switch_lp_equal_tmp_7_1 <= NMP_RunFSM_switch_lp_equal_tmp_21;
      while_while_nor_itm_2 <= while_while_nor_itm_1;
      NMP_RunFSM_switch_lp_equal_tmp_1_1 <= NMP_RunFSM_switch_lp_equal_tmp_22;
      NMP_RunFSM_switch_lp_equal_tmp_4_1 <= NMP_RunFSM_switch_lp_equal_tmp_23;
      NMP_RunFSM_switch_lp_equal_tmp_8_1 <= NMP_RunFSM_switch_lp_equal_tmp_24;
      NMP_RunFSM_switch_lp_equal_tmp_9_1 <= NMP_RunFSM_switch_lp_equal_tmp_25;
      NMP_RunFSM_switch_lp_equal_tmp_10_2 <= NMP_RunFSM_switch_lp_equal_tmp_10_1;
      NMP_RunFSM_switch_lp_equal_tmp_11_2 <= NMP_RunFSM_switch_lp_equal_tmp_11_1;
      NMP_RunFSM_switch_lp_equal_tmp_12_2 <= NMP_RunFSM_switch_lp_equal_tmp_12_1;
      NMP_RunFSM_switch_lp_or_tmp_1_1 <= NMP_RunFSM_switch_lp_or_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_config_vector_counter_sva <= 8'b00000000;
    end
    else if ( and_1063_tmp ) begin
      nmp_config_vector_counter_sva <= nmp_config_vector_counter_sva_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_config_num_vector_1_sva <= 8'b00000001;
      nmp_config_num_timestep_1_sva <= 16'b0000000000000001;
      nmp_config_mode_sva <= 3'b000;
      nmp_config_memory_index_1_sva <= 3'b000;
    end
    else if ( nmp_config_num_vector_1_and_cse ) begin
      nmp_config_num_vector_1_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[14:7];
      nmp_config_num_timestep_1_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[30:15];
      nmp_config_mode_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[3:1];
      nmp_config_memory_index_1_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[6:4];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_3_sva <= 1'b0;
      state_2_sva <= 1'b0;
      state_0_sva <= 1'b0;
      is_start_sva <= 1'b0;
    end
    else if ( state_and_cse ) begin
      state_3_sva <= next_state_3_lpi_1_dfm_4;
      state_2_sva <= next_state_2_lpi_1_dfm_4;
      state_0_sva <= next_state_0_lpi_1_dfm_4;
      is_start_sva <= NMP_RunFSM_switch_lp_mux_32_nl & (~ NMP_RunFSM_switch_lp_equal_tmp_10_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_1_sva <= 1'b0;
    end
    else if ( input_fixed_and_cse & nand_7_cse ) begin
      state_1_sva <= state_1_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_10_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_11_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_12_1 <= 1'b0;
      NMP_RunFSM_switch_lp_equal_tmp_1 <= 1'b0;
      nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1
          <= 1'b0;
      state_1_sva_dfm_1 <= 1'b0;
      while_while_nor_itm_1 <= 1'b0;
    end
    else if ( while_if_and_17_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= rva_in_PopNB_mioi_return_rsc_z_mxwt;
      NMP_RunFSM_switch_lp_equal_tmp_10_1 <= NMP_RunFSM_switch_lp_equal_tmp_13;
      NMP_RunFSM_switch_lp_equal_tmp_11_1 <= NMP_RunFSM_switch_lp_equal_tmp_14;
      NMP_RunFSM_switch_lp_equal_tmp_12_1 <= NMP_RunFSM_switch_lp_equal_tmp_15;
      NMP_RunFSM_switch_lp_equal_tmp_1 <= NMP_RunFSM_switch_lp_equal_tmp_16;
      nmp_config_UpdateVectorCounter_if_slc_nmp_config_UpdateVectorCounter_acc_9_1_svs_1
          <= operator_8_false_acc_1_itm_9_1;
      state_1_sva_dfm_1 <= MUX_s_1_2_2(next_state_1_lpi_1_dfm_4, state_1_sva_mx1,
          rva_in_PopNB_mioi_return_rsc_z_mxwt);
      while_while_nor_itm_1 <= (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) & rva_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_fixed_2_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_1_26_0_sva <= 27'b000000000000000000000000000;
      input_fixed_0_26_0_sva <= 27'b000000000000000000000000000;
    end
    else if ( and_1067_cse ) begin
      input_fixed_2_26_0_sva <= MUX_v_27_2_2(27'b000000000000000000000000000, NMP_ConvertInputToFixed_for_3_in_float_to_ac_fixed_lshift_1_itm,
          NMP_RunFSM_switch_lp_not_77_nl);
      input_fixed_1_26_0_sva <= MUX_v_27_2_2(27'b000000000000000000000000000, NMP_ConvertInputToFixed_for_2_in_float_to_ac_fixed_lshift_1_itm,
          NMP_RunFSM_switch_lp_not_78_nl);
      input_fixed_0_26_0_sva <= MUX_v_27_2_2(27'b000000000000000000000000000, NMP_ConvertInputToFixed_for_1_in_float_to_ac_fixed_lshift_1_itm,
          NMP_RunFSM_switch_lp_not_51_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_config_timestep_counter_sva <= 16'b0000000000000000;
    end
    else if ( and_1082_tmp ) begin
      nmp_config_timestep_counter_sva <= MUX_v_16_2_2(16'b0000000000000000, operator_16_false_acc_2_nl,
          mux_222_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_config_vector_counter_sva_3_1 <= 8'b00000000;
    end
    else if ( NMPRun_wen & (~ mux_tmp_6) & and_dcpl_172 & operator_8_false_acc_1_itm_9_1
        ) begin
      nmp_config_vector_counter_sva_3_1 <= nl_nmp_config_vector_counter_sva_3_1[7:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( NMPRun_wen & mux_cse & (~(NMP_RunFSM_switch_lp_equal_tmp_22 | NMP_RunFSM_switch_lp_equal_tmp_18_1
        | NMP_RunFSM_switch_lp_equal_tmp_20 | NMP_RunFSM_switch_lp_equal_tmp_23 |
        NMP_RunFSM_switch_lp_equal_tmp_17 | NMP_RunFSM_switch_lp_equal_tmp_19 | NMP_RunFSM_switch_lp_equal_tmp_21
        | NMP_RunFSM_switch_lp_equal_tmp_24 | NMP_RunFSM_switch_lp_equal_tmp_25 |
        NMP_RunFSM_switch_lp_equal_tmp_10_1 | NMP_RunFSM_switch_lp_equal_tmp_11_1
        | NMP_RunFSM_switch_lp_equal_tmp_12_1 | NMP_RunFSM_switch_lp_or_tmp_1)) &
        (~ or_dcpl_481) ) begin
      NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2 <= operator_3_false_operator_3_false_and_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_UpdateFSM_switch_lp_equal_tmp_1 <= 1'b0;
      NMP_UpdateFSM_switch_lp_equal_tmp_1_1 <= 1'b0;
      NMP_UpdateFSM_switch_lp_equal_tmp_4_1 <= 1'b0;
      NMP_UpdateFSM_switch_lp_or_tmp_1 <= 1'b0;
      NMP_UpdateFSM_switch_lp_nor_tmp_1 <= 1'b0;
      NMP_UpdateFSM_switch_lp_equal_tmp_2_1 <= 1'b0;
      NMP_UpdateFSM_switch_lp_equal_tmp_3_1 <= 1'b0;
      NMP_UpdateFSM_switch_lp_equal_tmp_5_1 <= 1'b0;
      NMP_UpdateFSM_switch_lp_equal_tmp_6_1 <= 1'b0;
    end
    else if ( NMP_UpdateFSM_switch_lp_and_4_cse ) begin
      NMP_UpdateFSM_switch_lp_equal_tmp_1 <= NMP_UpdateFSM_switch_lp_equal_tmp_7;
      NMP_UpdateFSM_switch_lp_equal_tmp_1_1 <= NMP_UpdateFSM_switch_lp_equal_tmp_8;
      NMP_UpdateFSM_switch_lp_equal_tmp_4_1 <= NMP_UpdateFSM_switch_lp_equal_tmp_9;
      NMP_UpdateFSM_switch_lp_or_tmp_1 <= NMP_UpdateFSM_switch_lp_or_tmp_1_1;
      NMP_UpdateFSM_switch_lp_nor_tmp_1 <= NMP_UpdateFSM_switch_lp_nor_tmp_1_1;
      NMP_UpdateFSM_switch_lp_equal_tmp_2_1 <= NMP_UpdateFSM_switch_lp_equal_tmp_10;
      NMP_UpdateFSM_switch_lp_equal_tmp_3_1 <= NMP_UpdateFSM_switch_lp_equal_tmp_11;
      NMP_UpdateFSM_switch_lp_equal_tmp_5_1 <= NMP_UpdateFSM_switch_lp_equal_tmp_12;
      NMP_UpdateFSM_switch_lp_equal_tmp_6_1 <= NMP_UpdateFSM_switch_lp_equal_tmp_13;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      next_state_3_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_481 | (~ fsm_output))) & (mux_tmp_6 | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
        | rva_in_PopNB_mioi_return_rsc_z_mxwt) ) begin
      next_state_3_lpi_1_dfm_3 <= next_state_3_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_itm_1
        | out_adp_set_value_ac_float_mux_80_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_2_itm_1
        | out_adp_set_value_ac_float_mux_81_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_3_itm_1
        | out_adp_set_value_ac_float_mux_82_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_4_itm_1
        | out_adp_set_value_ac_float_mux_83_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1
        | out_adp_set_value_ac_float_mux_84_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1
        | out_adp_set_value_ac_float_mux_85_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_7_itm_1
        | out_adp_set_value_ac_float_mux_86_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1
        | out_adp_set_value_ac_float_mux_87_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_9_itm_1
        | out_adp_set_value_ac_float_mux_88_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1
        | out_adp_set_value_ac_float_mux_89_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1
        | out_adp_set_value_ac_float_mux_90_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1
        | out_adp_set_value_ac_float_mux_91_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_13_itm_1
        | out_adp_set_value_ac_float_mux_92_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_14_itm_1
        | out_adp_set_value_ac_float_mux_93_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1
        | out_adp_set_value_ac_float_mux_94_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_483 | in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_16_itm_1
        | out_adp_set_value_ac_float_mux_95_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1
        | out_adp_set_value_ac_float_1_mux_80_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1
        | out_adp_set_value_ac_float_1_mux_81_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1
        | out_adp_set_value_ac_float_1_mux_82_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1
        | out_adp_set_value_ac_float_1_mux_83_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_5_itm_1
        | out_adp_set_value_ac_float_1_mux_84_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1
        | out_adp_set_value_ac_float_1_mux_85_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_7_itm_1
        | out_adp_set_value_ac_float_1_mux_86_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1
        | out_adp_set_value_ac_float_1_mux_87_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_9_itm_1
        | out_adp_set_value_ac_float_1_mux_88_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1
        | out_adp_set_value_ac_float_1_mux_89_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_11_itm_1
        | out_adp_set_value_ac_float_1_mux_90_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_12_itm_1
        | out_adp_set_value_ac_float_1_mux_91_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_13_itm_1
        | out_adp_set_value_ac_float_1_mux_92_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1
        | out_adp_set_value_ac_float_1_mux_93_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_15_itm_1
        | out_adp_set_value_ac_float_1_mux_94_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(or_dcpl_485 | or_dcpl_582 | in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_16_itm_1
        | out_adp_set_value_ac_float_1_mux_95_tmp_3)) ) begin
      NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs
          <= NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_3_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_16_tmp ) begin
      out_float_round_32_if_m_1_3_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_4_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_17_tmp ) begin
      out_float_round_32_if_m_1_4_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_5_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_18_tmp ) begin
      out_float_round_32_if_m_1_5_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_6_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_19_tmp ) begin
      out_float_round_32_if_m_1_6_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_7_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_20_tmp ) begin
      out_float_round_32_if_m_1_7_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_8_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_21_tmp ) begin
      out_float_round_32_if_m_1_8_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_9_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_22_tmp ) begin
      out_float_round_32_if_m_1_9_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_10_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_23_tmp ) begin
      out_float_round_32_if_m_1_10_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_11_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_24_tmp ) begin
      out_float_round_32_if_m_1_11_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_12_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_25_tmp ) begin
      out_float_round_32_if_m_1_12_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_13_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_26_tmp ) begin
      out_float_round_32_if_m_1_13_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_14_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_27_tmp ) begin
      out_float_round_32_if_m_1_14_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_15_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_28_tmp ) begin
      out_float_round_32_if_m_1_15_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_16_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_29_tmp ) begin
      out_float_round_32_if_m_1_16_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_17_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_30_tmp ) begin
      out_float_round_32_if_m_1_17_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_if_m_1_1_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_if_m_1_and_31_tmp ) begin
      out_float_round_32_if_m_1_1_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_3_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_16_tmp ) begin
      out_float_round_32_1_if_m_1_3_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_4_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_17_tmp ) begin
      out_float_round_32_1_if_m_1_4_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_5_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_18_tmp ) begin
      out_float_round_32_1_if_m_1_5_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_6_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_19_tmp ) begin
      out_float_round_32_1_if_m_1_6_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_7_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_20_tmp ) begin
      out_float_round_32_1_if_m_1_7_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_8_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_21_tmp ) begin
      out_float_round_32_1_if_m_1_8_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_9_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_22_tmp ) begin
      out_float_round_32_1_if_m_1_9_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_10_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_23_tmp ) begin
      out_float_round_32_1_if_m_1_10_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_11_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_24_tmp ) begin
      out_float_round_32_1_if_m_1_11_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_12_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_25_tmp ) begin
      out_float_round_32_1_if_m_1_12_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_13_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_26_tmp ) begin
      out_float_round_32_1_if_m_1_13_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_14_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_27_tmp ) begin
      out_float_round_32_1_if_m_1_14_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_15_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_28_tmp ) begin
      out_float_round_32_1_if_m_1_15_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_16_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_29_tmp ) begin
      out_float_round_32_1_if_m_1_16_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_17_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_30_tmp ) begin
      out_float_round_32_1_if_m_1_17_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_round_32_1_if_m_1_1_sva_1_3_0 <= 4'b0000;
    end
    else if ( out_float_round_32_1_if_m_1_and_31_tmp ) begin
      out_float_round_32_1_if_m_1_1_sva_1_3_0 <= NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_req_reg_write_data_data_6_4_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_6_4_sva_0 <= 1'b0;
      large_req_reg_write_data_data_14_12_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_14_12_sva_0 <= 1'b0;
      large_req_reg_write_data_data_22_20_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_22_20_sva_0 <= 1'b0;
      large_req_reg_write_data_data_30_28_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_30_28_sva_0 <= 1'b0;
      large_req_reg_write_data_data_38_36_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_38_36_sva_0 <= 1'b0;
      large_req_reg_write_data_data_46_44_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_46_44_sva_0 <= 1'b0;
      large_req_reg_write_data_data_54_52_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_54_52_sva_0 <= 1'b0;
      large_req_reg_write_data_data_62_60_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_62_60_sva_0 <= 1'b0;
      large_req_reg_write_data_data_70_68_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_70_68_sva_0 <= 1'b0;
      large_req_reg_write_data_data_78_76_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_78_76_sva_0 <= 1'b0;
      large_req_reg_write_data_data_86_84_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_86_84_sva_0 <= 1'b0;
      large_req_reg_write_data_data_94_92_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_94_92_sva_0 <= 1'b0;
      large_req_reg_write_data_data_102_100_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_102_100_sva_0 <= 1'b0;
      large_req_reg_write_data_data_110_108_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_110_108_sva_0 <= 1'b0;
      large_req_reg_write_data_data_118_116_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_118_116_sva_0 <= 1'b0;
      large_req_reg_write_data_data_126_124_sva_2_1 <= 2'b00;
      large_req_reg_write_data_data_126_124_sva_0 <= 1'b0;
    end
    else if ( large_req_reg_write_data_data_and_112_cse ) begin
      large_req_reg_write_data_data_6_4_sva_2_1 <= MUX_v_2_2_2(write_data_data_0_6_4_sva_dfm_1_2_1,
          write_data_data_0_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_6_4_sva_0 <= MUX_s_1_2_2(write_data_data_0_6_4_sva_dfm_1_0,
          write_data_data_0_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_14_12_sva_2_1 <= MUX_v_2_2_2(write_data_data_1_6_4_sva_dfm_1_2_1,
          write_data_data_1_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_14_12_sva_0 <= MUX_s_1_2_2(write_data_data_1_6_4_sva_dfm_1_0,
          write_data_data_1_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_22_20_sva_2_1 <= MUX_v_2_2_2(write_data_data_2_6_4_sva_dfm_1_2_1,
          write_data_data_2_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_22_20_sva_0 <= MUX_s_1_2_2(write_data_data_2_6_4_sva_dfm_1_0,
          write_data_data_2_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_30_28_sva_2_1 <= MUX_v_2_2_2(write_data_data_3_6_4_sva_dfm_1_2_1,
          write_data_data_3_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_30_28_sva_0 <= MUX_s_1_2_2(write_data_data_3_6_4_sva_dfm_1_0,
          write_data_data_3_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_38_36_sva_2_1 <= MUX_v_2_2_2(write_data_data_4_6_4_sva_dfm_1_2_1,
          write_data_data_4_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_38_36_sva_0 <= MUX_s_1_2_2(write_data_data_4_6_4_sva_dfm_1_0,
          write_data_data_4_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_46_44_sva_2_1 <= MUX_v_2_2_2(write_data_data_5_6_4_sva_dfm_1_2_1,
          write_data_data_5_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_46_44_sva_0 <= MUX_s_1_2_2(write_data_data_5_6_4_sva_dfm_1_0,
          write_data_data_5_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_54_52_sva_2_1 <= MUX_v_2_2_2(write_data_data_6_6_4_sva_dfm_1_2_1,
          write_data_data_6_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_54_52_sva_0 <= MUX_s_1_2_2(write_data_data_6_6_4_sva_dfm_1_0,
          write_data_data_6_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_62_60_sva_2_1 <= MUX_v_2_2_2(write_data_data_7_6_4_sva_dfm_1_2_1,
          write_data_data_7_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_62_60_sva_0 <= MUX_s_1_2_2(write_data_data_7_6_4_sva_dfm_1_0,
          write_data_data_7_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_70_68_sva_2_1 <= MUX_v_2_2_2(write_data_data_8_6_4_sva_dfm_1_2_1,
          write_data_data_8_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_70_68_sva_0 <= MUX_s_1_2_2(write_data_data_8_6_4_sva_dfm_1_0,
          write_data_data_8_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_78_76_sva_2_1 <= MUX_v_2_2_2(write_data_data_9_6_4_sva_dfm_1_2_1,
          write_data_data_9_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_78_76_sva_0 <= MUX_s_1_2_2(write_data_data_9_6_4_sva_dfm_1_0,
          write_data_data_9_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_86_84_sva_2_1 <= MUX_v_2_2_2(write_data_data_10_6_4_sva_dfm_1_2_1,
          write_data_data_10_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_86_84_sva_0 <= MUX_s_1_2_2(write_data_data_10_6_4_sva_dfm_1_0,
          write_data_data_10_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_94_92_sva_2_1 <= MUX_v_2_2_2(write_data_data_11_6_4_sva_dfm_1_2_1,
          write_data_data_11_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_94_92_sva_0 <= MUX_s_1_2_2(write_data_data_11_6_4_sva_dfm_1_0,
          write_data_data_11_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_102_100_sva_2_1 <= MUX_v_2_2_2(write_data_data_12_6_4_sva_dfm_1_2_1,
          write_data_data_12_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_102_100_sva_0 <= MUX_s_1_2_2(write_data_data_12_6_4_sva_dfm_1_0,
          write_data_data_12_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_110_108_sva_2_1 <= MUX_v_2_2_2(write_data_data_13_6_4_sva_dfm_1_2_1,
          write_data_data_13_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_110_108_sva_0 <= MUX_s_1_2_2(write_data_data_13_6_4_sva_dfm_1_0,
          write_data_data_13_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_118_116_sva_2_1 <= MUX_v_2_2_2(write_data_data_14_6_4_sva_dfm_1_2_1,
          write_data_data_14_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_118_116_sva_0 <= MUX_s_1_2_2(write_data_data_14_6_4_sva_dfm_1_0,
          write_data_data_14_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_126_124_sva_2_1 <= MUX_v_2_2_2(write_data_data_15_6_4_sva_dfm_1_2_1,
          write_data_data_15_6_4_sva_dfm_1_2_1_mx0w0, while_stage_0_19);
      large_req_reg_write_data_data_126_124_sva_0 <= MUX_s_1_2_2(write_data_data_15_6_4_sva_dfm_1_0,
          write_data_data_15_6_4_sva_dfm_1_0_mx0w0, while_stage_0_19);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      large_req_reg_write_data_data_7_sva <= 1'b0;
      large_req_reg_write_data_data_15_sva <= 1'b0;
      large_req_reg_write_data_data_23_sva <= 1'b0;
      large_req_reg_write_data_data_31_sva <= 1'b0;
      large_req_reg_write_data_data_39_sva <= 1'b0;
      large_req_reg_write_data_data_47_sva <= 1'b0;
      large_req_reg_write_data_data_55_sva <= 1'b0;
      large_req_reg_write_data_data_63_sva <= 1'b0;
      large_req_reg_write_data_data_71_sva <= 1'b0;
      large_req_reg_write_data_data_79_sva <= 1'b0;
      large_req_reg_write_data_data_87_sva <= 1'b0;
      large_req_reg_write_data_data_95_sva <= 1'b0;
      large_req_reg_write_data_data_103_sva <= 1'b0;
      large_req_reg_write_data_data_111_sva <= 1'b0;
      large_req_reg_write_data_data_119_sva <= 1'b0;
      large_req_reg_write_data_data_127_sva <= 1'b0;
    end
    else if ( large_req_reg_write_data_data_and_114_cse ) begin
      large_req_reg_write_data_data_7_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_860_mx0w0,
          write_data_data_0_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_15_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_863_mx0w0,
          write_data_data_1_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_23_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_866_mx0w0,
          write_data_data_2_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_31_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_869_mx0w0,
          write_data_data_3_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_39_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_872_mx0w0,
          write_data_data_4_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_47_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_875_mx0w0,
          write_data_data_5_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_55_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_878_mx0w0,
          write_data_data_6_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_63_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_881_mx0w0,
          write_data_data_7_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_71_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_884_mx0w0,
          write_data_data_8_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_79_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_887_mx0w0,
          write_data_data_9_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_87_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_890_mx0w0,
          write_data_data_10_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_95_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_893_mx0w0,
          write_data_data_11_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_103_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_896_mx0w0,
          write_data_data_12_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_111_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_899_mx0w0,
          write_data_data_13_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_119_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_902_mx0w0,
          write_data_data_14_7_sva_dfm_1, or_dcpl_471);
      large_req_reg_write_data_data_127_sva <= MUX_s_1_2_2(NMP_RunFSM_switch_lp_mux1h_905_mx0w0,
          write_data_data_15_7_sva_dfm_1, or_dcpl_471);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_1_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_15_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_1_sva_1 <= NMP_ConvertOutputToAdpfloat_for_1_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_2_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_14_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_2_sva_1 <= NMP_ConvertOutputToAdpfloat_for_2_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_3_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_13_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_3_sva_1 <= NMP_ConvertOutputToAdpfloat_for_3_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_4_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_12_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_4_sva_1 <= NMP_ConvertOutputToAdpfloat_for_4_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_5_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_11_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_5_sva_1 <= NMP_ConvertOutputToAdpfloat_for_5_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_6_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_10_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_6_sva_1 <= NMP_ConvertOutputToAdpfloat_for_6_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_7_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_9_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_7_sva_1 <= NMP_ConvertOutputToAdpfloat_for_7_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_8_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_8_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_8_sva_1 <= NMP_ConvertOutputToAdpfloat_for_8_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_9_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_7_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_9_sva_1 <= NMP_ConvertOutputToAdpfloat_for_9_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_10_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_6_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_10_sva_1 <= NMP_ConvertOutputToAdpfloat_for_10_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_11_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_5_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_11_sva_1 <= NMP_ConvertOutputToAdpfloat_for_11_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_12_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_4_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_12_sva_1 <= NMP_ConvertOutputToAdpfloat_for_12_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_13_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_3_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_13_sva_1 <= NMP_ConvertOutputToAdpfloat_for_13_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_14_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_2_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_14_sva_1 <= NMP_ConvertOutputToAdpfloat_for_14_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_15_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_1_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_15_sva_1 <= NMP_ConvertOutputToAdpfloat_for_15_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_215 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_less_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_sva_1 <= NMP_ConvertOutputToAdpfloat_for_16_leading_sign_32_1_1_0_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_1_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_15_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_1_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_1_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_2_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_14_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_2_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_2_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_3_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_13_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_3_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_3_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_4_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_12_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_4_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_4_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_5_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_11_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_5_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_5_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_6_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_10_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_6_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_6_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_7_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_9_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_7_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_7_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_8_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_8_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_8_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_8_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_9_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_7_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_9_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_9_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_10_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_6_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_10_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_10_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_11_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_5_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_11_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_11_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_12_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_4_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_12_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_12_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_13_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_3_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_13_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_13_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_14_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_2_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_14_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_14_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_15_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_1_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_15_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_15_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_sva_1 <= 5'b00000;
    end
    else if ( NMPRun_wen & and_dcpl_217 & and_dcpl_249 & out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_less_tmp
        ) begin
      out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_sva_1 <= NMP_ConvertOutputToAdpfloat_1_for_16_leading_sign_32_1_1_0_2_out_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_psp_sva
          <= 11'b00000000000;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_5_enex5
        ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_psp_sva
          <= nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_psp_sva[10:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_9_0
          <= 10'b0000000000;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_6_enex5
        ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_9_0
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_mx0w0[9:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TR000000
          <= 10'b0000000000;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5
        ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TR000000
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_itm
          <= 11'b00000000000;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_5_enex5
        ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_itm
          <= nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_itm[10:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4 <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp )
        begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4 <= MUX1HOT_v_7_5_2(ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_3,
          7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, {(~ NMP_RunFSM_switch_lp_conc_itm_7_1)
          , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_cse , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_1_cse
          , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_2_cse , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_3_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      max_value_26_0_sva_26 <= 1'b0;
    end
    else if ( while_if_and_12_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      max_value_26_0_sva_26 <= NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_54_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      max_value_26_0_sva_25_0 <= 26'b00000000000000000000000000;
    end
    else if ( and_1085_enex5 & (~ or_924_itm) ) begin
      max_value_26_0_sva_25_0 <= NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_52_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_cse <= 27'b000000000000000000000000000;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_cse <= NMP_ComputeSoftmaxExp_for_asn_30_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      max_value_26_0_sva_dfm_13_1_26 <= 1'b0;
    end
    else if ( max_value_and_1_cse ) begin
      max_value_26_0_sva_dfm_13_1_26 <= MUX_s_1_2_2(max_value_26_0_sva_dfm_12_26_mx0,
          (NMP_ComputeSoftmaxExp_for_asn_28_itm_2[26]), NMP_ComputeSoftmaxMax_for_if_less_2_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxMax_for_asn_13_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 ) begin
      NMP_ComputeSoftmaxMax_for_asn_13_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_29_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      max_value_26_0_sva_dfm_13_1_25_0 <= 26'b00000000000000000000000000;
    end
    else if ( max_value_and_enex5 ) begin
      max_value_26_0_sva_dfm_13_1_25_0 <= MUX_v_26_2_2(max_value_26_0_sva_dfm_12_25_0_mx0,
          (NMP_ComputeSoftmaxExp_for_asn_28_itm_2[25:0]), NMP_ComputeSoftmaxMax_for_if_less_2_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_30_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_66_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_30_itm_2 <= NMP_RunFSM_switch_lp_asn_104_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_29_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_67_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_29_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_29_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_28_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_68_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_28_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_28_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_27_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_69_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_27_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_27_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_26_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_70_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_26_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_26_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_25_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_21_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_25_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_25_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_24_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_71_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_24_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_24_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_23_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_72_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_23_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_23_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_22_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_73_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_22_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_22_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_21_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_74_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_21_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_21_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_20_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_75_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_20_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_20_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_19_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_76_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_19_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_19_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_18_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_77_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_18_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_18_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_17_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_78_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_17_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_17_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_16_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_79_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_16_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_16_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_80_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_config_is_valid_sva <= 1'b0;
    end
    else if ( NMPRun_wen & (~(nmp_config_ConfigRead_unequal_tmp_1 | or_dcpl_694 |
        nand_7_cse | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt))) ) begin
      nmp_config_is_valid_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nmp_config_adpbias_1_ftd <= 1'b0;
      reg_nmp_config_adpbias_1_ftd_1 <= 2'b00;
    end
    else if ( nmp_config_adpbias_1_and_ssc ) begin
      reg_nmp_config_adpbias_1_ftd <= nmp_config_adpbias_1_sva_dfm_3_1_2;
      reg_nmp_config_adpbias_1_ftd_1 <= MUX_v_2_2_2(nmp_config_adpbias_1_sva_dfm_3_1_1_0,
          (nmp_config_memory_index_1_sva[1:0]), and_671_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      next_state_1_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( NMPRun_wen & (~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | rva_in_PopNB_mioi_return_rsc_z_mxwt))
        ) begin
      next_state_1_lpi_1_dfm_3 <= next_state_1_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_16 <= 1'b0;
    end
    else if ( NMPRun_wen & while_stage_0_17 & (~ while_while_nor_itm_15) ) begin
      while_while_and_itm_16 <= while_while_and_itm_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      sum_exp_39_4_sva_st_1 <= 36'b000000000000000000000000000000000000;
    end
    else if ( sum_exp_and_3_enex5 ) begin
      sum_exp_39_4_sva_st_1 <= sum_exp_39_4_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_0_3_itm_3
          <= 1'b0;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_6_cse )
        begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_0_3_itm_3
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_0_3_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_16 <= 2'b00;
      NMP_PrepareWriteReq_asn_1_itm_15_rsp_0 <= 1'b0;
      reg_NMP_PrepareWriteReq_asn_1_itm_15_1_ftd <= 1'b0;
    end
    else if ( NMP_PrepareWriteReq_and_15_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_16 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_15;
      NMP_PrepareWriteReq_asn_1_itm_15_rsp_0 <= NMP_PrepareWriteReq_asn_1_itm_14_7;
      reg_NMP_PrepareWriteReq_asn_1_itm_15_1_ftd <= NMP_PrepareWriteReq_asn_1_itm_14_6_0_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_45_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_96_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_45_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_45_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_43_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_97_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_43_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_43_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_41_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_98_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_41_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_41_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_39_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_99_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_39_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_39_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_37_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_100_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_37_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_37_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_35_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_101_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_35_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_35_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_33_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_102_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_33_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_33_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_31_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_103_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_31_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_31_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_29_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_104_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_29_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_29_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_27_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_105_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_27_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_27_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_25_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_106_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_25_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_25_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_23_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_107_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_23_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_23_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_21_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_108_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_21_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_21_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_19_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_109_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_19_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_19_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_17_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_110_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_17_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_17_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_itm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_111_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_itm_3 <= NMP_ComputeSoftmaxNormalize_for_asn_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_2 <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_2_enex5
        ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_2 <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_161_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_9 <= NMP_ComputeRMSNormalize_for_asn_60_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_162_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_9 <= NMP_ComputeRMSNormalize_for_asn_58_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_163_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_9 <= NMP_ComputeRMSNormalize_for_asn_56_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_164_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_9 <= NMP_ComputeRMSNormalize_for_asn_54_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_165_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_9 <= NMP_ComputeRMSNormalize_for_asn_52_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_166_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_9 <= NMP_ComputeRMSNormalize_for_asn_50_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_167_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_9 <= NMP_ComputeRMSNormalize_for_asn_48_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_168_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_9 <= NMP_ComputeRMSNormalize_for_asn_46_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_169_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_9 <= NMP_ComputeRMSNormalize_for_asn_44_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_170_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_9 <= NMP_ComputeRMSNormalize_for_asn_42_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_171_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_9 <= NMP_ComputeRMSNormalize_for_asn_40_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_172_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_9 <= NMP_ComputeRMSNormalize_for_asn_38_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_173_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_9 <= NMP_ComputeRMSNormalize_for_asn_36_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_174_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_10 <= NMP_ComputeRMSNormalize_for_asn_34_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_175_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_10 <= NMP_ComputeRMSNormalize_for_asn_32_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_10 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_176_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_10 <= NMP_ComputeRMSNormalize_for_asn_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_2
          <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_4_enex5
        ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_2
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_16 <= 2'b00;
      reg_NMP_PrepareReadReq_asn_2_itm_15_ftd_1 <= 3'b000;
      NMP_PrepareReadReq_asn_1_itm_15_7_6_rsp_0 <= 1'b0;
      NMP_PrepareReadReq_asn_1_itm_15_7_6_rsp_1 <= 1'b0;
    end
    else if ( NMP_PrepareReadReq_and_17_cse ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_16 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_15;
      reg_NMP_PrepareReadReq_asn_2_itm_15_ftd_1 <= NMP_PrepareReadReq_asn_2_itm_14_15_7_rsp_1;
      NMP_PrepareReadReq_asn_1_itm_15_7_6_rsp_0 <= reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_1_1;
      NMP_PrepareReadReq_asn_1_itm_15_7_6_rsp_1 <= reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_16 <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_16_ftd <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_16_ftd_1 <= 2'b00;
      rva_out_reg_data_10_8_sva_dfm_3_16 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_16 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_12_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_16 <= rva_out_reg_data_0_sva_dfm_3_15;
      reg_rva_out_reg_data_98_96_sva_dfm_3_16_ftd <= rva_out_reg_data_98_96_sva_dfm_3_15_rsp_0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_16_ftd_1 <= rva_out_reg_data_98_96_sva_dfm_3_15_rsp_1;
      rva_out_reg_data_10_8_sva_dfm_3_16 <= rva_out_reg_data_10_8_sva_dfm_3_15;
      rva_out_reg_data_34_32_sva_dfm_3_16 <= rva_out_reg_data_34_32_sva_dfm_3_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_16 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_104_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_16 <= rva_out_reg_data_79_64_sva_dfm_3_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_16 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_105_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_16 <= rva_out_reg_data_55_48_sva_dfm_3_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_3
          <= 1'b0;
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_4
          <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_129_cse ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_3
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_2_1;
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_4
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_3_39
          <= 1'b0;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_2_cse
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_3_39
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_2_39;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= 1'b0;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse ) begin
      NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_sva_1 | (NMP_ConvertOutputToAdpfloat_for_16_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_15_sva_1 | (NMP_ConvertOutputToAdpfloat_for_15_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_14_sva_1 | (NMP_ConvertOutputToAdpfloat_for_14_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_13_sva_1 | (NMP_ConvertOutputToAdpfloat_for_13_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_12_sva_1 | (NMP_ConvertOutputToAdpfloat_for_12_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_11_sva_1 | (NMP_ConvertOutputToAdpfloat_for_11_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_10_sva_1 | (NMP_ConvertOutputToAdpfloat_for_10_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_9_sva_1 | (NMP_ConvertOutputToAdpfloat_for_9_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_8_sva_1 | (NMP_ConvertOutputToAdpfloat_for_8_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_7_sva_1 | (NMP_ConvertOutputToAdpfloat_for_7_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_6_sva_1 | (NMP_ConvertOutputToAdpfloat_for_6_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_5_sva_1 | (NMP_ConvertOutputToAdpfloat_for_5_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_4_sva_1 | (NMP_ConvertOutputToAdpfloat_for_4_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_3_sva_1 | (NMP_ConvertOutputToAdpfloat_for_3_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_2_sva_1 | (NMP_ConvertOutputToAdpfloat_for_2_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs
          <= (NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_for_out_float_m_4_1_sva_1 | (NMP_ConvertOutputToAdpfloat_for_1_out_float_round_32_if_m_1_acc_tmp[3:0]!=4'b0000)));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
      NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= 1'b0;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse ) begin
      NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_16_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_15_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_15_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_14_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_14_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_13_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_13_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_12_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_12_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_11_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_11_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_10_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_10_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_9_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_9_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_8_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_8_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_7_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_7_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_6_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_6_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_5_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_5_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_4_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_4_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_3_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_3_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_2_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_2_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
      NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs
          <= (NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp[6])
          & (~(NMP_ConvertOutputToAdpfloat_1_for_out_float_m_4_1_sva_1 | (NMP_ConvertOutputToAdpfloat_1_for_1_out_float_round_32_1_if_m_1_acc_tmp[3:0]!=4'b0000)));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_itm
          <= 10'b0000000000;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_itm
          <= 10'b0000000000;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_itm
          <= 8'b00000000;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_1_cse
        ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_itm
          <= z_out_1;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_itm
          <= z_out_2[35:26];
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_itm
          <= z_out;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_itm
          <= 10'b0000000000;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_itm
          <= 10'b0000000000;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_itm
          <= 8'b00000000;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_2_cse
        ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_itm
          <= z_out_1;
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_itm
          <= z_out_2[35:26];
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_itm
          <= z_out;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      sum_exp_39_4_sva_3_34_0 <= 35'b00000000000000000000000000000000000;
    end
    else if ( sum_exp_and_4_enex5 ) begin
      sum_exp_39_4_sva_3_34_0 <= sum_exp_39_4_sva_2[34:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxSum_for_acc_7_itm_1 <= 34'b0000000000000000000000000000000000;
      NMP_ComputeSoftmaxSum_for_acc_8_itm_1 <= 34'b0000000000000000000000000000000000;
      NMP_ComputeSoftmaxSum_for_acc_9_itm_1 <= 34'b0000000000000000000000000000000000;
      NMP_ComputeSoftmaxSum_for_acc_11_itm_1 <= 34'b0000000000000000000000000000000000;
      NMP_ComputeSoftmaxSum_for_acc_12_itm_1 <= 33'b000000000000000000000000000000000;
      NMP_ComputeSoftmaxSum_for_acc_13_itm_1 <= 33'b000000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxSum_for_and_cse ) begin
      NMP_ComputeSoftmaxSum_for_acc_7_itm_1 <= nl_NMP_ComputeSoftmaxSum_for_acc_7_itm_1[33:0];
      NMP_ComputeSoftmaxSum_for_acc_8_itm_1 <= nl_NMP_ComputeSoftmaxSum_for_acc_8_itm_1[33:0];
      NMP_ComputeSoftmaxSum_for_acc_9_itm_1 <= nl_NMP_ComputeSoftmaxSum_for_acc_9_itm_1[33:0];
      NMP_ComputeSoftmaxSum_for_acc_11_itm_1 <= nl_NMP_ComputeSoftmaxSum_for_acc_11_itm_1[33:0];
      NMP_ComputeSoftmaxSum_for_acc_12_itm_1 <= nl_NMP_ComputeSoftmaxSum_for_acc_12_itm_1[32:0];
      NMP_ComputeSoftmaxSum_for_acc_13_itm_1 <= nl_NMP_ComputeSoftmaxSum_for_acc_13_itm_1[32:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1
          <= 20'b00000000000000000000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_8_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1
          <= ({ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_11_8
          , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_7_6
          , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_5_0})
          * ({2'b10 , NMP_PrepareWriteReq_asn_1_itm_5_5_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mux_1_itm_2
          <= 10'b0000000000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_9_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mux_1_itm_2
          <= NMP_PrepareReadReq_asn_2_itm_5_9_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      max_value_26_0_sva_dfm_9_1_26 <= 1'b0;
    end
    else if ( max_value_and_3_cse ) begin
      max_value_26_0_sva_dfm_9_1_26 <= max_value_26_0_sva_dfm_9_1_26_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxMax_for_if_less_5_itm_1 <= 1'b0;
    end
    else if ( NMP_ComputeSoftmaxMax_for_if_and_tmp ) begin
      NMP_ComputeSoftmaxMax_for_if_less_5_itm_1 <= NMP_ComputeSoftmaxMax_for_if_less_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      max_value_26_0_sva_dfm_9_1_25_0 <= 26'b00000000000000000000000000;
    end
    else if ( max_value_and_9_enex5 ) begin
      max_value_26_0_sva_dfm_9_1_25_0 <= max_value_26_0_sva_dfm_9_1_25_0_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nmp_config_adpbias_1_sva_dfm_3_1_2 <= 1'b0;
      nmp_config_adpbias_1_sva_dfm_3_1_1_0 <= 2'b00;
    end
    else if ( nmp_config_adpbias_1_and_1_ssc ) begin
      nmp_config_adpbias_1_sva_dfm_3_1_2 <= MUX1HOT_s_1_3_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[33]),
          nmp_config_adpbias_1_sva_mx1_2, rva_out_reg_data_98_96_sva_dfm_3_1_2, {nmp_config_adpbias_1_sva_dfm_3_1_mx0c0
          , nmp_config_adpbias_1_sva_dfm_3_1_mx0c1 , nmp_config_adpbias_1_sva_dfm_3_1_mx0c2});
      nmp_config_adpbias_1_sva_dfm_3_1_1_0 <= MUX1HOT_v_2_3_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[32:31]),
          nmp_config_adpbias_1_sva_mx1_1_0, rva_out_reg_data_98_96_sva_dfm_3_1_1_0,
          {nmp_config_adpbias_1_sva_dfm_3_1_mx0c0 , nmp_config_adpbias_1_sva_dfm_3_1_mx0c1
          , nmp_config_adpbias_1_sva_dfm_3_1_mx0c2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_15 <= 1'b0;
    end
    else if ( NMPRun_wen & while_stage_0_16 & (~ while_while_nor_itm_14) ) begin
      while_while_and_itm_15 <= while_while_and_itm_14;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_0_3_itm_2
          <= 1'b0;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_7_cse )
        begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_slc_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_0_3_itm_2
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_15 <= 2'b00;
      NMP_PrepareWriteReq_asn_1_itm_14_7 <= 1'b0;
      NMP_PrepareWriteReq_asn_1_itm_14_6_0_rsp_0 <= 1'b0;
    end
    else if ( NMP_PrepareWriteReq_and_18_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_15 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_14;
      NMP_PrepareWriteReq_asn_1_itm_14_7 <= reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd;
      NMP_PrepareWriteReq_asn_1_itm_14_6_0_rsp_0 <= reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd_1_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_45_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_112_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_45_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_45_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_43_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_113_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_43_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_43_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_41_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_114_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_41_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_41_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_39_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_115_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_39_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_39_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_37_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_116_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_37_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_37_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_35_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_117_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_35_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_35_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_33_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_118_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_33_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_33_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_31_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_119_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_31_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_31_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_29_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_120_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_29_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_29_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_27_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_121_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_27_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_27_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_25_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_122_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_25_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_25_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_23_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_123_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_23_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_23_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_21_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_124_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_21_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_21_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_19_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_125_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_19_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_19_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_17_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_126_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_17_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_17_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_itm_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_127_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_itm_2 <= NMP_ComputeSoftmaxNormalize_for_asn_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_29_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_81_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_29_itm_1 <= input_fixed_14_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_28_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_82_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_28_itm_1 <= input_fixed_13_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_27_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_83_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_27_itm_1 <= input_fixed_12_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_26_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_84_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_26_itm_1 <= input_fixed_11_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_25_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_85_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_25_itm_1 <= input_fixed_10_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_24_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_86_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_24_itm_1 <= input_fixed_9_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_23_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_87_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_23_itm_1 <= input_fixed_8_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_22_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_88_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_22_itm_1 <= input_fixed_7_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_21_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_89_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_21_itm_1 <= input_fixed_6_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_20_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_90_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_20_itm_1 <= input_fixed_5_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_19_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_91_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_19_itm_1 <= input_fixed_4_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_18_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_92_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_18_itm_1 <= input_fixed_3_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_17_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_93_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_17_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_17_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_16_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_94_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_16_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_16_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_itm_2 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_95_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_itm_2 <= NMP_ComputeSoftmaxExp_for_asn_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_177_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_8 <= NMP_ComputeRMSNormalize_for_asn_60_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_178_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_8 <= NMP_ComputeRMSNormalize_for_asn_58_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_179_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_8 <= NMP_ComputeRMSNormalize_for_asn_56_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_180_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_8 <= NMP_ComputeRMSNormalize_for_asn_54_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_181_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_8 <= NMP_ComputeRMSNormalize_for_asn_52_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_182_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_8 <= NMP_ComputeRMSNormalize_for_asn_50_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_183_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_8 <= NMP_ComputeRMSNormalize_for_asn_48_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_184_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_8 <= NMP_ComputeRMSNormalize_for_asn_46_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_185_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_8 <= NMP_ComputeRMSNormalize_for_asn_44_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_186_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_8 <= NMP_ComputeRMSNormalize_for_asn_42_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_187_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_8 <= NMP_ComputeRMSNormalize_for_asn_40_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_188_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_8 <= NMP_ComputeRMSNormalize_for_asn_38_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_189_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_8 <= NMP_ComputeRMSNormalize_for_asn_36_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_190_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_9 <= NMP_ComputeRMSNormalize_for_asn_34_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_191_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_9 <= NMP_ComputeRMSNormalize_for_asn_32_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_9 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_192_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_9 <= NMP_ComputeRMSNormalize_for_asn_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_1 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_56_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_1 <= NMP_PrepareReadReq_asn_1_itm_13_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_15 <= 2'b00;
      reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_1_1 <= 1'b0;
      reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_0 <= 1'b0;
      NMP_PrepareReadReq_asn_2_itm_14_15_7_rsp_1 <= 3'b000;
    end
    else if ( NMP_PrepareReadReq_and_20_cse ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_15 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_14;
      reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_1_1 <= reg_NMP_PrepareReadReq_asn_1_itm_13_ftd;
      reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_0 <= reg_NMP_PrepareReadReq_asn_1_itm_13_ftd_1;
      NMP_PrepareReadReq_asn_2_itm_14_15_7_rsp_1 <= reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_15 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_15 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_15 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_15_rsp_0 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_15_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_18_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_15 <= rva_out_reg_data_0_sva_dfm_3_14;
      rva_out_reg_data_10_8_sva_dfm_3_15 <= rva_out_reg_data_10_8_sva_dfm_3_14;
      rva_out_reg_data_34_32_sva_dfm_3_15 <= rva_out_reg_data_34_32_sva_dfm_3_14;
      rva_out_reg_data_98_96_sva_dfm_3_15_rsp_0 <= rva_out_reg_data_98_96_sva_dfm_3_14_2;
      rva_out_reg_data_98_96_sva_dfm_3_15_rsp_1 <= rva_out_reg_data_98_96_sva_dfm_3_14_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_15 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_106_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_15 <= rva_out_reg_data_79_64_sva_dfm_3_14;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_15 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_107_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_15 <= rva_out_reg_data_55_48_sva_dfm_3_14;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_2_1
          <= 1'b0;
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_3
          <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_135_cse ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_2_1
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_1;
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_3
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_3 <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_13_enex5
        ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_3 <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_2_39
          <= 1'b0;
    end
    else if ( NMPRun_wen & and_dcpl_137 & and_dcpl_134 & (~ NMP_RunFSM_switch_lp_equal_tmp_10)
        & NMP_RunFSM_switch_lp_equal_tmp_3_9 & ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_1
        & (~ NMP_RunFSM_switch_lp_conc_itm_10_0) ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_2_39
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_1_39;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm
          <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_cse )
        begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm
          <= MUX_v_7_2_2(7'b0000000, ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_qif_acc_cse,
          ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_or_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      operator_40_0_false_AC_TRN_AC_WRAP_1_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_38_0_itm
          <= 39'b000000000000000000000000000000000000000;
    end
    else if ( operator_40_0_false_AC_TRN_AC_WRAP_1_and_enex5 ) begin
      operator_40_0_false_AC_TRN_AC_WRAP_1_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_38_0_itm
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_38_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_tmp
        ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_qif_acc_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      sum_exp_39_4_sva_2 <= 36'b000000000000000000000000000000000000;
    end
    else if ( sum_exp_and_5_enex5 ) begin
      sum_exp_39_4_sva_2 <= sum_exp_39_4_sva_st_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      exp_values_15_sva <= 32'b00000000000000000000000000000000;
      exp_values_14_sva <= 32'b00000000000000000000000000000000;
      exp_values_13_sva <= 32'b00000000000000000000000000000000;
      exp_values_12_sva <= 32'b00000000000000000000000000000000;
      exp_values_11_sva <= 32'b00000000000000000000000000000000;
      exp_values_10_sva <= 32'b00000000000000000000000000000000;
      exp_values_9_sva <= 32'b00000000000000000000000000000000;
      exp_values_8_sva <= 32'b00000000000000000000000000000000;
      exp_values_7_sva <= 32'b00000000000000000000000000000000;
      exp_values_6_sva <= 32'b00000000000000000000000000000000;
      exp_values_5_sva <= 32'b00000000000000000000000000000000;
      exp_values_4_sva <= 32'b00000000000000000000000000000000;
      exp_values_3_sva <= 32'b00000000000000000000000000000000;
      exp_values_2_sva <= 32'b00000000000000000000000000000000;
      exp_values_1_sva <= 32'b00000000000000000000000000000000;
      exp_values_0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( and_1094_cse ) begin
      exp_values_15_sva <= exp_values_15_sva_mx1;
      exp_values_14_sva <= exp_values_14_sva_mx1;
      exp_values_13_sva <= exp_values_13_sva_mx1;
      exp_values_12_sva <= exp_values_12_sva_mx1;
      exp_values_11_sva <= exp_values_11_sva_mx1;
      exp_values_10_sva <= exp_values_10_sva_mx1;
      exp_values_9_sva <= exp_values_9_sva_mx1;
      exp_values_8_sva <= exp_values_8_sva_mx1;
      exp_values_7_sva <= exp_values_7_sva_mx1;
      exp_values_6_sva <= exp_values_6_sva_mx1;
      exp_values_5_sva <= exp_values_5_sva_mx1;
      exp_values_4_sva <= exp_values_4_sva_mx1;
      exp_values_3_sva <= exp_values_3_sva_mx1;
      exp_values_2_sva <= exp_values_2_sva_mx1;
      exp_values_1_sva <= exp_values_1_sva_mx1;
      exp_values_0_sva <= exp_values_0_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_62_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_63_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_16_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_2_itm_1
          <= 3'b000;
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_58_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_59_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_15_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_6_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_7_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_2_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_54_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_55_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_14_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_3_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_50_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_51_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_13_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_4_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_46_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_47_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_12_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_18_itm_1
          <= 3'b000;
      NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_5_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_42_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_43_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_11_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_22_itm_1
          <= 3'b000;
      NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_6_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_38_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_39_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_26_itm_1
          <= 3'b000;
      NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_7_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_34_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_35_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_9_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
      NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= 9'b000000000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_30_itm_1
          <= 3'b000;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_31_itm_1
          <= 7'b0000000;
      NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= 10'b0000000000;
      NMP_ComputeSoftmaxExp_for_8_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= 9'b000000000;
    end
    else if ( ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_9_cse
        ) begin
      NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_62_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_63_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z[33:32]);
      NMP_ComputeSoftmaxExp_for_16_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_16_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z[42:34];
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_1_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_2_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[33:32]);
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_1_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[42:34];
      NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_15_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_58_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_59_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z[33:32]);
      NMP_ComputeSoftmaxExp_for_15_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_15_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_15_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z[42:34];
      NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_2_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_6_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_7_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z[33:32]);
      NMP_ComputeSoftmaxExp_for_2_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_2_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_2_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z[42:34];
      NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_14_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_54_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_55_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z[33:32]);
      NMP_ComputeSoftmaxExp_for_14_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_14_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_14_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z[42:34];
      NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_3_sva_1[18:10];
      NMP_ComputeSoftmaxExp_for_3_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_3_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_3_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z[42:34];
      NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_13_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_50_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_51_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z[33:32]);
      NMP_ComputeSoftmaxExp_for_13_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_13_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_13_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z[42:34];
      NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_4_sva_1[18:10];
      NMP_ComputeSoftmaxExp_for_4_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_4_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_4_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[42:34];
      NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_12_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_46_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_47_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z[33:32]);
      NMP_ComputeSoftmaxExp_for_12_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_12_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_12_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z[42:34];
      NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_5_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_18_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[33:32]);
      NMP_ComputeSoftmaxExp_for_5_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_5_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_5_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[42:34];
      NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_11_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_42_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_43_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z[33:32]);
      NMP_ComputeSoftmaxExp_for_11_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_11_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_11_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z[42:34];
      NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_6_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_22_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[33:32]);
      NMP_ComputeSoftmaxExp_for_6_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_6_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_6_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z[42:34];
      NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_10_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_38_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_39_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z[33:32]);
      NMP_ComputeSoftmaxExp_for_10_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_10_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_7_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_26_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[33:32]);
      NMP_ComputeSoftmaxExp_for_7_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_7_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_7_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[42:34];
      NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_34_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_35_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z[33:32]);
      NMP_ComputeSoftmaxExp_for_9_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_9_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z[42:34];
      NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000000
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_8_sva_1[18:10];
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_30_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z[33:32]);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_31_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z[33:32]);
      NMP_ComputeSoftmaxExp_for_8_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_000001
          <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mul_psp_8_sva_1[9:0];
      NMP_ComputeSoftmaxExp_for_8_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_input_inter_32_8_24_12_itm_1
          <= NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z[42:34];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      max_value_26_0_sva_dfm_6_1_26 <= 1'b0;
      max_value_26_0_sva_dfm_6_1_25_0 <= 26'b00000000000000000000000000;
    end
    else if ( max_value_and_5_cse ) begin
      max_value_26_0_sva_dfm_6_1_26 <= MUX_s_1_2_2(max_value_26_0_sva_dfm_5_26_mx0,
          (input_fixed_6_26_0_sva[26]), NMP_ComputeSoftmaxMax_for_if_less_9_itm);
      max_value_26_0_sva_dfm_6_1_25_0 <= MUX_v_26_2_2(max_value_26_0_sva_dfm_5_25_0_mx0,
          (input_fixed_6_26_0_sva[25:0]), NMP_ComputeSoftmaxMax_for_if_less_9_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_14 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ while_while_nor_itm_13) & while_stage_0_15 ) begin
      while_while_and_itm_14 <= while_while_and_itm_13;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_RunFSM_switch_lp_asn_104_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_RunFSM_switch_lp_and_342_enex5 ) begin
      NMP_RunFSM_switch_lp_asn_104_itm_1 <= input_fixed_15_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_13_ftd <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_63_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_13_ftd <= NMP_PrepareWriteReq_asn_2_itm_12_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_13_ftd_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareWriteReq_and_64_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_13_ftd_1 <= NMP_PrepareWriteReq_asn_2_itm_12_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd <= 1'b0;
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_14 <= 2'b00;
      reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd_1_6 <= 1'b0;
    end
    else if ( NMP_PrepareWriteReq_and_21_cse ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd <= NMP_PrepareWriteReq_asn_1_itm_12_rsp_0;
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_14 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_13;
      reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd_1_6 <= reg_NMP_PrepareWriteReq_asn_1_itm_12_1_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_adp_set_value_ac_float_1_asn_15_itm_13_ftd <= 1'b0;
      reg_out_adp_set_value_ac_float_1_asn_15_itm_13_ftd_1 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_3_ssc ) begin
      reg_out_adp_set_value_ac_float_1_asn_15_itm_13_ftd <= out_adp_set_value_ac_float_1_asn_15_itm_12_rsp_0;
      reg_out_adp_set_value_ac_float_1_asn_15_itm_13_ftd_1 <= out_adp_set_value_ac_float_1_asn_15_itm_12_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_45_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_128_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_45_itm_1 <= exp_values_15_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_43_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_129_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_43_itm_1 <= exp_values_14_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_41_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_130_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_41_itm_1 <= exp_values_13_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_39_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_131_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_39_itm_1 <= exp_values_12_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_37_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_132_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_37_itm_1 <= exp_values_11_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_35_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_133_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_35_itm_1 <= exp_values_10_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_33_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_134_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_33_itm_1 <= exp_values_9_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_31_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_135_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_31_itm_1 <= exp_values_8_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_29_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_136_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_29_itm_1 <= exp_values_7_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_27_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_137_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_27_itm_1 <= exp_values_6_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_25_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_138_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_25_itm_1 <= exp_values_5_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_23_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_139_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_23_itm_1 <= exp_values_4_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_21_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_140_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_21_itm_1 <= exp_values_3_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_19_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_141_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_19_itm_1 <= exp_values_2_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_17_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_142_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_17_itm_1 <= exp_values_1_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_143_enex5 ) begin
      NMP_ComputeSoftmaxNormalize_for_asn_itm_1 <= exp_values_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_17_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_96_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_17_itm_1 <= input_fixed_2_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_16_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_97_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_16_itm_1 <= input_fixed_1_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxExp_for_asn_itm_1 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_98_enex5 ) begin
      NMP_ComputeSoftmaxExp_for_asn_itm_1 <= input_fixed_0_26_0_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_13_ftd <= 1'b0;
      reg_out_adp_set_value_ac_float_asn_15_itm_13_ftd_1 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_and_3_ssc ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_13_ftd <= out_adp_set_value_ac_float_asn_15_itm_12_rsp_0;
      reg_out_adp_set_value_ac_float_asn_15_itm_13_ftd_1 <= out_adp_set_value_ac_float_asn_15_itm_12_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_193_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_7 <= NMP_ComputeRMSNormalize_for_asn_60_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_194_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_7 <= NMP_ComputeRMSNormalize_for_asn_58_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_195_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_7 <= NMP_ComputeRMSNormalize_for_asn_56_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_196_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_7 <= NMP_ComputeRMSNormalize_for_asn_54_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_197_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_7 <= NMP_ComputeRMSNormalize_for_asn_52_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_198_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_7 <= NMP_ComputeRMSNormalize_for_asn_50_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_199_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_7 <= NMP_ComputeRMSNormalize_for_asn_48_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_200_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_7 <= NMP_ComputeRMSNormalize_for_asn_46_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_201_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_7 <= NMP_ComputeRMSNormalize_for_asn_44_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_202_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_7 <= NMP_ComputeRMSNormalize_for_asn_42_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_203_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_7 <= NMP_ComputeRMSNormalize_for_asn_40_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_204_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_7 <= NMP_ComputeRMSNormalize_for_asn_38_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_205_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_7 <= NMP_ComputeRMSNormalize_for_asn_36_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_206_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_8 <= NMP_ComputeRMSNormalize_for_asn_34_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_207_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_8 <= NMP_ComputeRMSNormalize_for_asn_32_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_8 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_208_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_8 <= NMP_ComputeRMSNormalize_for_asn_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareReadReq_and_57_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_1 <= NMP_PrepareReadReq_asn_2_itm_12_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_14 <= 2'b00;
      reg_NMP_PrepareReadReq_asn_1_itm_13_ftd <= 1'b0;
      reg_NMP_PrepareReadReq_asn_1_itm_13_ftd_1 <= 1'b0;
      reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_2_0 <= 3'b000;
    end
    else if ( NMP_PrepareReadReq_and_23_cse ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_14 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_13;
      reg_NMP_PrepareReadReq_asn_1_itm_13_ftd <= NMP_PrepareReadReq_asn_1_itm_12_7_6_rsp_0;
      reg_NMP_PrepareReadReq_asn_1_itm_13_ftd_1 <= NMP_PrepareReadReq_asn_1_itm_12_7_6_rsp_1;
      reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_2_0 <= reg_NMP_PrepareReadReq_asn_2_itm_12_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_14 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_14 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_14 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_14_2 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_14_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_24_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_14 <= rva_out_reg_data_0_sva_dfm_3_13;
      rva_out_reg_data_10_8_sva_dfm_3_14 <= rva_out_reg_data_10_8_sva_dfm_3_13;
      rva_out_reg_data_34_32_sva_dfm_3_14 <= rva_out_reg_data_34_32_sva_dfm_3_13;
      rva_out_reg_data_98_96_sva_dfm_3_14_2 <= reg_rva_out_reg_data_98_96_sva_dfm_3_13_ftd;
      rva_out_reg_data_98_96_sva_dfm_3_14_1_0 <= reg_rva_out_reg_data_98_96_sva_dfm_3_13_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_14 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_108_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_14 <= rva_out_reg_data_79_64_sva_dfm_3_13;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_14 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_109_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_14 <= rva_out_reg_data_55_48_sva_dfm_3_13;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_1
          <= 1'b0;
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_2
          <= 1'b0;
    end
    else if ( NMP_RunFSM_switch_lp_and_158_cse ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_1
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_2;
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_2
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_2 <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_14_enex5
        ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_2 <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_1_39
          <= 1'b0;
    end
    else if ( NMPRun_wen & and_dcpl_145 & ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_or_tmp_2
        & (~ NMP_RunFSM_switch_lp_equal_tmp_9) & NMP_RunFSM_switch_lp_equal_tmp_3_8
        & NMP_RunFSM_switch_lp_conc_itm_9_2 & (~ NMP_RunFSM_switch_lp_conc_itm_9_3)
        & (~(NMP_RunFSM_switch_lp_conc_itm_9_1 | NMP_RunFSM_switch_lp_conc_itm_9_0))
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_1_39
          <= operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp[39];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_or_itm
          <= 1'b0;
    end
    else if ( NMPRun_wen & (~(((operator_40_16_false_AC_TRN_AC_WRAP_lshift_tmp==40'b0000000000000000000000000000000000000000))
        | (~ while_stage_0_11) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
        | (~ NMP_RunFSM_switch_lp_conc_itm_9_2) | NMP_RunFSM_switch_lp_conc_itm_9_3
        | NMP_RunFSM_switch_lp_conc_itm_9_1 | NMP_RunFSM_switch_lp_conc_itm_9_0))
        ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_or_itm
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_mx0_39
          | (ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_mx0_38_0!=39'b000000000000000000000000000000000000000);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      max_value_26_0_sva_dfm_2_1_26 <= 1'b0;
    end
    else if ( max_value_and_7_cse ) begin
      max_value_26_0_sva_dfm_2_1_26 <= max_value_26_0_sva_dfm_2_1_26_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeSoftmaxMax_for_if_less_12_itm_1 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ state_0_sva) & state_2_sva & (~ state_3_sva) & and_dcpl_443
        ) begin
      NMP_ComputeSoftmaxMax_for_if_less_12_itm_1 <= NMP_ComputeSoftmaxMax_for_if_less_12_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      max_value_26_0_sva_dfm_2_1_25_0 <= 26'b00000000000000000000000000;
    end
    else if ( max_value_and_10_enex5 ) begin
      max_value_26_0_sva_dfm_2_1_25_0 <= max_value_26_0_sva_dfm_2_1_25_0_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_13 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ while_while_nor_itm_12) & while_stage_0_14 ) begin
      while_while_and_itm_13 <= while_while_and_itm_12;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_13 <= 2'b00;
      NMP_PrepareWriteReq_asn_1_itm_12_rsp_0 <= 1'b0;
      reg_NMP_PrepareWriteReq_asn_1_itm_12_1_ftd <= 1'b0;
    end
    else if ( NMP_PrepareWriteReq_and_24_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_13 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_12;
      NMP_PrepareWriteReq_asn_1_itm_12_rsp_0 <= NMP_PrepareWriteReq_asn_1_itm_11_7;
      reg_NMP_PrepareWriteReq_asn_1_itm_12_1_ftd <= NMP_PrepareWriteReq_asn_1_itm_11_6_0_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_209_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_6 <= NMP_ComputeRMSNormalize_for_asn_60_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_210_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_6 <= NMP_ComputeRMSNormalize_for_asn_58_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_211_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_6 <= NMP_ComputeRMSNormalize_for_asn_56_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_212_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_6 <= NMP_ComputeRMSNormalize_for_asn_54_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_213_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_6 <= NMP_ComputeRMSNormalize_for_asn_52_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_214_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_6 <= NMP_ComputeRMSNormalize_for_asn_50_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_215_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_6 <= NMP_ComputeRMSNormalize_for_asn_48_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_216_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_6 <= NMP_ComputeRMSNormalize_for_asn_46_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_217_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_6 <= NMP_ComputeRMSNormalize_for_asn_44_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_218_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_6 <= NMP_ComputeRMSNormalize_for_asn_42_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_219_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_6 <= NMP_ComputeRMSNormalize_for_asn_40_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_220_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_6 <= NMP_ComputeRMSNormalize_for_asn_38_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_221_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_6 <= NMP_ComputeRMSNormalize_for_asn_36_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_222_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_7 <= NMP_ComputeRMSNormalize_for_asn_34_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_223_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_7 <= NMP_ComputeRMSNormalize_for_asn_32_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_7 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_224_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_7 <= NMP_ComputeRMSNormalize_for_asn_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_13 <= 2'b00;
      reg_NMP_PrepareReadReq_asn_2_itm_12_ftd_1 <= 3'b000;
      NMP_PrepareReadReq_asn_1_itm_12_7_6_rsp_0 <= 1'b0;
      NMP_PrepareReadReq_asn_1_itm_12_7_6_rsp_1 <= 1'b0;
    end
    else if ( NMP_PrepareReadReq_and_26_cse ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_13 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_12;
      reg_NMP_PrepareReadReq_asn_2_itm_12_ftd_1 <= NMP_PrepareReadReq_asn_2_itm_11_15_7_rsp_1;
      NMP_PrepareReadReq_asn_1_itm_12_7_6_rsp_0 <= NMP_PrepareReadReq_asn_1_itm_11_7;
      NMP_PrepareReadReq_asn_1_itm_12_7_6_rsp_1 <= NMP_PrepareReadReq_asn_1_itm_11_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_13 <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_13_ftd <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_13_ftd_1 <= 2'b00;
      rva_out_reg_data_10_8_sva_dfm_3_13 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_13 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_30_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_13 <= rva_out_reg_data_0_sva_dfm_3_12;
      reg_rva_out_reg_data_98_96_sva_dfm_3_13_ftd <= rva_out_reg_data_98_96_sva_dfm_3_12_rsp_0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_13_ftd_1 <= rva_out_reg_data_98_96_sva_dfm_3_12_rsp_1;
      rva_out_reg_data_10_8_sva_dfm_3_13 <= rva_out_reg_data_10_8_sva_dfm_3_12;
      rva_out_reg_data_34_32_sva_dfm_3_13 <= rva_out_reg_data_34_32_sva_dfm_3_12;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_13 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_110_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_13 <= rva_out_reg_data_79_64_sva_dfm_3_12;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_13 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_111_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_13 <= rva_out_reg_data_55_48_sva_dfm_3_12;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_1
          <= 1'b0;
    end
    else if ( NMPRun_wen & and_dcpl_154 & (~ NMP_RunFSM_switch_lp_equal_tmp_8) )
        begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_or_tmp_1
          <= (sum_exp_39_4_sva_1!=36'b000000000000000000000000000000000000);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1 <= 7'b0000000;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_9_cse )
        begin
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1 <= nl_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1[6:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      sum_sq_1_39_4_sva <= 36'b000000000000000000000000000000000000;
    end
    else if ( (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_3
        | (~ while_stage_0_5) | (~(NMP_RunFSM_switch_lp_equal_tmp_3 | NMP_RunFSM_switch_lp_equal_tmp_2_2)))
        & (NMP_RunFSM_switch_lp_equal_tmp_2_3 | NMP_RunFSM_switch_lp_equal_tmp_4)
        & input_fixed_and_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 ) begin
      sum_sq_1_39_4_sva <= sum_sq_1_39_4_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      sum_sq_1_39_4_sva_2_1 <= 36'b000000000000000000000000000000000000;
    end
    else if ( NMPRun_wen & and_dcpl_169 & NMP_RunFSM_switch_lp_equal_tmp_2_2 & (~
        NMP_RunFSM_switch_lp_equal_tmp_3) ) begin
      sum_sq_1_39_4_sva_2_1 <= readslicef_40_36_4(NMP_ComputeRMSSumSq_for_acc_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_12 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ while_while_nor_itm_11) & while_stage_0_13 ) begin
      while_while_and_itm_12 <= while_while_and_itm_11;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_12 <= 2'b00;
      NMP_PrepareWriteReq_asn_1_itm_11_7 <= 1'b0;
      NMP_PrepareWriteReq_asn_1_itm_11_6_0_rsp_0 <= 1'b0;
    end
    else if ( NMP_PrepareWriteReq_and_27_ssc ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_12 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_11;
      NMP_PrepareWriteReq_asn_1_itm_11_7 <= reg_NMP_PrepareWriteReq_asn_1_itm_10_ftd;
      NMP_PrepareWriteReq_asn_1_itm_11_6_0_rsp_0 <= reg_NMP_PrepareWriteReq_asn_1_itm_10_1_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_225_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_5 <= NMP_ComputeRMSNormalize_for_asn_60_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_226_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_5 <= NMP_ComputeRMSNormalize_for_asn_58_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_227_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_5 <= NMP_ComputeRMSNormalize_for_asn_56_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_228_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_5 <= NMP_ComputeRMSNormalize_for_asn_54_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_229_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_5 <= NMP_ComputeRMSNormalize_for_asn_52_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_230_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_5 <= NMP_ComputeRMSNormalize_for_asn_50_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_231_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_5 <= NMP_ComputeRMSNormalize_for_asn_48_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_232_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_5 <= NMP_ComputeRMSNormalize_for_asn_46_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_233_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_5 <= NMP_ComputeRMSNormalize_for_asn_44_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_234_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_5 <= NMP_ComputeRMSNormalize_for_asn_42_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_235_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_5 <= NMP_ComputeRMSNormalize_for_asn_40_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_236_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_5 <= NMP_ComputeRMSNormalize_for_asn_38_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_237_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_5 <= NMP_ComputeRMSNormalize_for_asn_36_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_238_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_6 <= NMP_ComputeRMSNormalize_for_asn_34_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_239_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_6 <= NMP_ComputeRMSNormalize_for_asn_32_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_6 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_240_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_6 <= NMP_ComputeRMSNormalize_for_asn_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_12 <= 2'b00;
      NMP_PrepareReadReq_asn_1_itm_11_7 <= 1'b0;
      NMP_PrepareReadReq_asn_1_itm_11_6 <= 1'b0;
      NMP_PrepareReadReq_asn_2_itm_11_15_7_rsp_1 <= 3'b000;
    end
    else if ( NMP_PrepareReadReq_and_29_ssc ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_12 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_11;
      NMP_PrepareReadReq_asn_1_itm_11_7 <= reg_NMP_PrepareReadReq_asn_1_itm_10_ftd;
      NMP_PrepareReadReq_asn_1_itm_11_6 <= reg_NMP_PrepareReadReq_asn_1_itm_10_ftd_1;
      NMP_PrepareReadReq_asn_2_itm_11_15_7_rsp_1 <= reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_12 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_12 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_12 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_12_rsp_0 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_12_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_36_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_12 <= rva_out_reg_data_0_sva_dfm_3_11;
      rva_out_reg_data_10_8_sva_dfm_3_12 <= rva_out_reg_data_10_8_sva_dfm_3_11;
      rva_out_reg_data_34_32_sva_dfm_3_12 <= rva_out_reg_data_34_32_sva_dfm_3_11;
      rva_out_reg_data_98_96_sva_dfm_3_12_rsp_0 <= rva_out_reg_data_98_96_sva_dfm_3_11_2;
      rva_out_reg_data_98_96_sva_dfm_3_12_rsp_1 <= rva_out_reg_data_98_96_sva_dfm_3_11_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_12 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_112_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_12 <= rva_out_reg_data_79_64_sva_dfm_3_11;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_12 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_113_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_12 <= rva_out_reg_data_55_48_sva_dfm_3_11;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_11 <= 1'b0;
    end
    else if ( NMPRun_wen & while_stage_0_12 & (~ while_while_nor_itm_10) ) begin
      while_while_and_itm_11 <= while_while_and_itm_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_10_ftd <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_65_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_10_ftd <= NMP_PrepareWriteReq_asn_2_itm_9_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_10_ftd_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareWriteReq_and_66_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_10_ftd_1 <= NMP_PrepareWriteReq_asn_2_itm_9_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_10_ftd <= 1'b0;
      reg_NMP_PrepareWriteReq_asn_1_itm_10_1_ftd <= 1'b0;
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_11 <= 2'b00;
    end
    else if ( NMP_PrepareWriteReq_and_30_ssc ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_10_ftd <= NMP_PrepareWriteReq_asn_1_itm_9_rsp_0;
      reg_NMP_PrepareWriteReq_asn_1_itm_10_1_ftd <= NMP_PrepareWriteReq_asn_1_itm_9_rsp_1_rsp_0;
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_11 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_10_1_ftd_1 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_67_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_10_1_ftd_1 <= NMP_PrepareWriteReq_asn_1_itm_9_rsp_1_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_adp_set_value_ac_float_1_asn_15_itm_10_ftd <= 1'b0;
      reg_out_adp_set_value_ac_float_1_asn_15_itm_10_ftd_1 <= 2'b00;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_32_cse ) begin
      reg_out_adp_set_value_ac_float_1_asn_15_itm_10_ftd <= out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_0;
      reg_out_adp_set_value_ac_float_1_asn_15_itm_10_ftd_1 <= out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_10_ftd <= 1'b0;
      reg_out_adp_set_value_ac_float_asn_15_itm_10_ftd_1 <= 2'b00;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_32_cse ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_10_ftd <= out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_0;
      reg_out_adp_set_value_ac_float_asn_15_itm_10_ftd_1 <= out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_241_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_60_itm_4 <= reg_NMP_RunFSM_switch_lp_asn_104_itm_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_242_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_4 <= NMP_ComputeRMSNormalize_for_asn_58_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_243_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_4 <= NMP_ComputeRMSNormalize_for_asn_56_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_244_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_4 <= NMP_ComputeRMSNormalize_for_asn_54_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_245_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_4 <= NMP_ComputeRMSNormalize_for_asn_52_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_246_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_4 <= NMP_ComputeRMSNormalize_for_asn_50_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_247_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_4 <= NMP_ComputeRMSNormalize_for_asn_48_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_248_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_4 <= NMP_ComputeRMSNormalize_for_asn_46_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_249_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_4 <= NMP_ComputeRMSNormalize_for_asn_44_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_250_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_4 <= NMP_ComputeRMSNormalize_for_asn_42_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_251_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_4 <= NMP_ComputeRMSNormalize_for_asn_40_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_252_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_4 <= NMP_ComputeRMSNormalize_for_asn_38_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_253_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_4 <= NMP_ComputeRMSNormalize_for_asn_36_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_254_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_5 <= NMP_ComputeRMSNormalize_for_asn_34_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_255_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_5 <= NMP_ComputeRMSNormalize_for_asn_32_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_5 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_256_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_5 <= NMP_ComputeRMSNormalize_for_asn_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_2 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_58_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_2 <= NMP_PrepareReadReq_asn_2_itm_9_rsp_0_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_3 <= 3'b000;
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_11 <= 2'b00;
    end
    else if ( NMP_PrepareReadReq_and_32_ssc ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_3 <= NMP_PrepareReadReq_asn_2_itm_9_rsp_0_rsp_1;
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_11 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareReadReq_and_59_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_1 <= NMP_PrepareReadReq_asn_2_itm_9_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_11 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_11 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_11 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_11_2 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_11_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_42_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_11 <= rva_out_reg_data_0_sva_dfm_3_10;
      rva_out_reg_data_10_8_sva_dfm_3_11 <= rva_out_reg_data_10_8_sva_dfm_3_10;
      rva_out_reg_data_34_32_sva_dfm_3_11 <= rva_out_reg_data_34_32_sva_dfm_3_10;
      rva_out_reg_data_98_96_sva_dfm_3_11_2 <= reg_rva_out_reg_data_98_96_sva_dfm_3_10_ftd;
      rva_out_reg_data_98_96_sva_dfm_3_11_1_0 <= reg_rva_out_reg_data_98_96_sva_dfm_3_10_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_11 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_114_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_11 <= rva_out_reg_data_79_64_sva_dfm_3_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_11 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_115_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_11 <= rva_out_reg_data_55_48_sva_dfm_3_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_10 <= 1'b0;
    end
    else if ( NMPRun_wen & while_stage_0_11 & (~ while_while_nor_itm_9) ) begin
      while_while_and_itm_10 <= while_while_and_itm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_10 <= 2'b00;
      NMP_PrepareWriteReq_asn_1_itm_9_rsp_0 <= 1'b0;
      NMP_PrepareWriteReq_asn_1_itm_9_rsp_1_rsp_0 <= 1'b0;
    end
    else if ( NMP_PrepareWriteReq_and_35_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_10 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_9;
      NMP_PrepareWriteReq_asn_1_itm_9_rsp_0 <= NMP_PrepareWriteReq_asn_1_itm_8_7;
      NMP_PrepareWriteReq_asn_1_itm_9_rsp_1_rsp_0 <= NMP_PrepareWriteReq_asn_1_itm_8_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_257_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_58_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_29_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_258_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_56_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_28_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_259_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_54_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_27_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_260_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_52_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_26_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_261_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_50_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_25_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_262_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_48_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_24_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_263_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_46_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_23_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_264_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_44_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_22_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_265_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_42_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_21_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_266_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_40_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_20_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_267_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_38_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_19_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_268_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_36_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_18_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_269_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_4 <= NMP_ComputeRMSNormalize_for_asn_34_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_270_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_32_itm_4 <= NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_26_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_4 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_271_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_4 <= NMP_ComputeRMSNormalize_for_asn_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_10 <= 2'b00;
      NMP_PrepareReadReq_asn_1_itm_9_rsp_0 <= 1'b0;
      NMP_PrepareReadReq_asn_2_itm_9_rsp_0_rsp_1 <= 3'b000;
      NMP_PrepareReadReq_asn_1_itm_9_rsp_1_rsp_0 <= 1'b0;
    end
    else if ( NMP_PrepareReadReq_and_36_cse ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_10 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_9;
      NMP_PrepareReadReq_asn_1_itm_9_rsp_0 <= NMP_PrepareReadReq_asn_1_itm_8_7;
      NMP_PrepareReadReq_asn_2_itm_9_rsp_0_rsp_1 <= NMP_PrepareReadReq_asn_2_itm_8_9_7;
      NMP_PrepareReadReq_asn_1_itm_9_rsp_1_rsp_0 <= NMP_PrepareReadReq_asn_1_itm_8_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_10 <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_10_ftd <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_10_ftd_1 <= 2'b00;
      rva_out_reg_data_10_8_sva_dfm_3_10 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_10 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_48_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_10 <= rva_out_reg_data_0_sva_dfm_3_9;
      reg_rva_out_reg_data_98_96_sva_dfm_3_10_ftd <= rva_out_reg_data_98_96_sva_dfm_3_9_rsp_0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_10_ftd_1 <= rva_out_reg_data_98_96_sva_dfm_3_9_rsp_1;
      rva_out_reg_data_10_8_sva_dfm_3_10 <= rva_out_reg_data_10_8_sva_dfm_3_9;
      rva_out_reg_data_34_32_sva_dfm_3_10 <= rva_out_reg_data_34_32_sva_dfm_3_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_10 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_116_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_10 <= rva_out_reg_data_79_64_sva_dfm_3_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_10 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_117_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_10 <= rva_out_reg_data_55_48_sva_dfm_3_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_9 <= 1'b0;
    end
    else if ( NMPRun_wen & while_stage_0_10 & (~ while_while_nor_itm_8) ) begin
      while_while_and_itm_9 <= while_while_and_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_9 <= 2'b00;
      NMP_PrepareWriteReq_asn_1_itm_8_7 <= 1'b0;
      NMP_PrepareWriteReq_asn_1_itm_8_6 <= 1'b0;
    end
    else if ( NMP_PrepareWriteReq_and_38_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_9 <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_14_itm_1_1_0;
      NMP_PrepareWriteReq_asn_1_itm_8_7 <= NMP_PrepareWriteReq_asn_1_itm_7_7;
      NMP_PrepareWriteReq_asn_1_itm_8_6 <= NMP_PrepareWriteReq_asn_1_itm_7_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_272_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_34_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_17_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_3 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_273_enex5 ) begin
      NMP_ComputeRMSNormalize_for_asn_itm_3 <= NMP_ComputeSoftmaxExp_for_asn_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_9 <= 2'b00;
      NMP_PrepareReadReq_asn_1_itm_8_7 <= 1'b0;
      NMP_PrepareReadReq_asn_2_itm_8_9_7 <= 3'b000;
      NMP_PrepareReadReq_asn_1_itm_8_6 <= 1'b0;
    end
    else if ( NMP_PrepareReadReq_and_39_cse ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_9 <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_1_0;
      NMP_PrepareReadReq_asn_1_itm_8_7 <= NMP_PrepareReadReq_asn_1_itm_7_7;
      NMP_PrepareReadReq_asn_2_itm_8_9_7 <= reg_NMP_PrepareReadReq_asn_2_itm_7_ftd_1;
      NMP_PrepareReadReq_asn_1_itm_8_6 <= NMP_PrepareReadReq_asn_1_itm_7_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_9 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_9 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_9 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_9_rsp_0 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_9_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_54_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_9 <= rva_out_reg_data_0_sva_dfm_3_8;
      rva_out_reg_data_10_8_sva_dfm_3_9 <= rva_out_reg_data_10_8_sva_dfm_3_8;
      rva_out_reg_data_34_32_sva_dfm_3_9 <= rva_out_reg_data_34_32_sva_dfm_3_8;
      rva_out_reg_data_98_96_sva_dfm_3_9_rsp_0 <= rva_out_reg_data_98_96_sva_dfm_3_8_2;
      rva_out_reg_data_98_96_sva_dfm_3_9_rsp_1 <= rva_out_reg_data_98_96_sva_dfm_3_8_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_9 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_118_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_9 <= rva_out_reg_data_79_64_sva_dfm_3_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_9 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_119_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_9 <= rva_out_reg_data_55_48_sva_dfm_3_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_8 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ while_while_nor_itm_7) & while_stage_0_9 ) begin
      while_while_and_itm_8 <= while_while_and_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_8 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_8 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_8 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_8_2 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_8_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_60_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_8 <= rva_out_reg_data_0_sva_dfm_3_7;
      rva_out_reg_data_10_8_sva_dfm_3_8 <= rva_out_reg_data_10_8_sva_dfm_3_7;
      rva_out_reg_data_34_32_sva_dfm_3_8 <= rva_out_reg_data_34_32_sva_dfm_3_7;
      rva_out_reg_data_98_96_sva_dfm_3_8_2 <= reg_rva_out_reg_data_98_96_sva_dfm_3_7_ftd;
      rva_out_reg_data_98_96_sva_dfm_3_8_1_0 <= reg_rva_out_reg_data_98_96_sva_dfm_3_7_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_8 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_120_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_8 <= rva_out_reg_data_79_64_sva_dfm_3_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_8 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_121_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_8 <= rva_out_reg_data_55_48_sva_dfm_3_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_7 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ while_while_nor_itm_6) & while_stage_0_8 ) begin
      while_while_and_itm_7 <= while_while_and_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_6 <= 16'b0000000000000000;
    end
    else if ( NMP_PrepareWriteReq_and_68_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_6 <= NMP_PrepareWriteReq_asn_2_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_7 <= 2'b00;
      NMP_PrepareWriteReq_asn_1_itm_6_7_6 <= 2'b00;
    end
    else if ( NMP_PrepareWriteReq_and_41_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_7 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_6;
      NMP_PrepareWriteReq_asn_1_itm_6_7_6 <= NMP_PrepareWriteReq_asn_1_itm_5_7_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_7 <= 2'b00;
      NMP_PrepareReadReq_asn_1_itm_6_rsp_0 <= 2'b00;
    end
    else if ( NMP_PrepareReadReq_and_44_cse ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_7 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_6;
      NMP_PrepareReadReq_asn_1_itm_6_rsp_0 <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_7_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_7 <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_7_ftd <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_7_ftd_1 <= 2'b00;
      rva_out_reg_data_10_8_sva_dfm_3_7 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_7 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_66_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_7 <= rva_out_reg_data_0_sva_dfm_3_6;
      reg_rva_out_reg_data_98_96_sva_dfm_3_7_ftd <= rva_out_reg_data_98_96_sva_dfm_3_6_rsp_0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_7_ftd_1 <= rva_out_reg_data_98_96_sva_dfm_3_6_rsp_1;
      rva_out_reg_data_10_8_sva_dfm_3_7 <= rva_out_reg_data_10_8_sva_dfm_3_6;
      rva_out_reg_data_34_32_sva_dfm_3_7 <= rva_out_reg_data_34_32_sva_dfm_3_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_7 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_122_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_7 <= rva_out_reg_data_79_64_sva_dfm_3_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_7 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_123_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_7 <= rva_out_reg_data_55_48_sva_dfm_3_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_6 <= 1'b0;
    end
    else if ( NMPRun_wen & while_stage_0_7 & (~ while_while_nor_itm_5) ) begin
      while_while_and_itm_6 <= while_while_and_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_5 <= 16'b0000000000000000;
    end
    else if ( NMP_PrepareWriteReq_and_69_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_5 <= NMP_PrepareWriteReq_asn_2_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_6 <= 2'b00;
    end
    else if ( NMP_PrepareWriteReq_and_44_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_6 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_6 <= 2'b00;
    end
    else if ( NMPRun_wen & and_dcpl_354 & and_dcpl_482 & (~ NMP_RunFSM_switch_lp_conc_itm_5_2)
        ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_6 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_6 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_6 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_6 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_6_rsp_0 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_6_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_72_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_6 <= rva_out_reg_data_0_sva_dfm_3_5;
      rva_out_reg_data_10_8_sva_dfm_3_6 <= rva_out_reg_data_10_8_sva_dfm_3_5;
      rva_out_reg_data_34_32_sva_dfm_3_6 <= rva_out_reg_data_34_32_sva_dfm_3_5;
      rva_out_reg_data_98_96_sva_dfm_3_6_rsp_0 <= rva_out_reg_data_98_96_sva_dfm_3_5_2;
      rva_out_reg_data_98_96_sva_dfm_3_6_rsp_1 <= rva_out_reg_data_98_96_sva_dfm_3_5_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_124_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_6 <= rva_out_reg_data_79_64_sva_dfm_3_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_6 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_125_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_6 <= rva_out_reg_data_55_48_sva_dfm_3_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_5 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ while_while_nor_itm_4) & while_stage_0_6 ) begin
      while_while_and_itm_5 <= while_while_and_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_4 <= 16'b0000000000000000;
    end
    else if ( NMP_PrepareWriteReq_and_70_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_4 <= NMP_PrepareWriteReq_asn_2_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_4 <= 8'b00000000;
    end
    else if ( NMP_PrepareWriteReq_and_71_enex5 ) begin
      NMP_PrepareWriteReq_asn_1_itm_4 <= NMP_PrepareWriteReq_asn_1_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_5 <= 2'b00;
    end
    else if ( NMP_PrepareWriteReq_and_47_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_5 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_adp_set_value_ac_float_1_asn_15_itm_4_ftd <= 1'b0;
      reg_out_adp_set_value_ac_float_1_asn_15_itm_4_ftd_1 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_11_ssc ) begin
      reg_out_adp_set_value_ac_float_1_asn_15_itm_4_ftd <= out_adp_set_value_ac_float_1_asn_15_itm_3_rsp_0;
      reg_out_adp_set_value_ac_float_1_asn_15_itm_4_ftd_1 <= out_adp_set_value_ac_float_1_asn_15_itm_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_4_ftd <= 1'b0;
      reg_out_adp_set_value_ac_float_asn_15_itm_4_ftd_1 <= 2'b00;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_128_cse ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_4_ftd <= out_adp_set_value_ac_float_asn_15_itm_3_rsp_0;
      reg_out_adp_set_value_ac_float_asn_15_itm_4_ftd_1 <= out_adp_set_value_ac_float_asn_15_itm_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_4 <= 16'b0000000000000000;
    end
    else if ( NMP_PrepareReadReq_and_60_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_4 <= NMP_PrepareReadReq_asn_2_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_5 <= 2'b00;
    end
    else if ( NMP_PrepareReadReq_and_47_cse ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_5 <= NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_5 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_5 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_5 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_5_2 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_5_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_78_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_5 <= rva_out_reg_data_0_sva_dfm_3_4;
      rva_out_reg_data_10_8_sva_dfm_3_5 <= rva_out_reg_data_10_8_sva_dfm_3_4;
      rva_out_reg_data_34_32_sva_dfm_3_5 <= rva_out_reg_data_34_32_sva_dfm_3_4;
      rva_out_reg_data_98_96_sva_dfm_3_5_2 <= reg_rva_out_reg_data_98_96_sva_dfm_3_4_ftd;
      rva_out_reg_data_98_96_sva_dfm_3_5_1_0 <= reg_rva_out_reg_data_98_96_sva_dfm_3_4_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_126_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_5 <= rva_out_reg_data_79_64_sva_dfm_3_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_5 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_127_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_5 <= rva_out_reg_data_55_48_sva_dfm_3_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_4 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ while_while_nor_itm_3) & while_stage_0_5 ) begin
      while_while_and_itm_4 <= while_while_and_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_3 <= 16'b0000000000000000;
    end
    else if ( NMP_PrepareWriteReq_and_72_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_3 <= NMP_PrepareWriteReq_asn_2_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_3 <= 8'b00000000;
    end
    else if ( NMP_PrepareWriteReq_and_73_enex5 ) begin
      NMP_PrepareWriteReq_asn_1_itm_3 <= NMP_PrepareWriteReq_asn_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_4 <= 2'b00;
    end
    else if ( NMP_PrepareWriteReq_and_50_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_4 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_3 <= 16'b0000000000000000;
    end
    else if ( NMP_PrepareReadReq_and_61_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_3 <= NMP_PrepareWriteReq_asn_2_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_3 <= 8'b00000000;
    end
    else if ( NMP_PrepareReadReq_and_62_enex5 ) begin
      NMP_PrepareReadReq_asn_1_itm_3 <= NMP_PrepareWriteReq_asn_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_4 <= 2'b00;
    end
    else if ( NMP_PrepareReadReq_and_50_cse ) begin
      NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_4 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_4 <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_4_ftd <= 1'b0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_4_ftd_1 <= 2'b00;
      rva_out_reg_data_10_8_sva_dfm_3_4 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_4 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_84_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_4 <= rva_out_reg_data_0_sva_dfm_3_3;
      reg_rva_out_reg_data_98_96_sva_dfm_3_4_ftd <= rva_out_reg_data_98_96_sva_dfm_3_3_rsp_0;
      reg_rva_out_reg_data_98_96_sva_dfm_3_4_ftd_1 <= rva_out_reg_data_98_96_sva_dfm_3_3_rsp_1;
      rva_out_reg_data_10_8_sva_dfm_3_4 <= rva_out_reg_data_10_8_sva_dfm_3_3;
      rva_out_reg_data_34_32_sva_dfm_3_4 <= rva_out_reg_data_34_32_sva_dfm_3_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_128_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_4 <= rva_out_reg_data_79_64_sva_dfm_3_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_129_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_4 <= rva_out_reg_data_55_48_sva_dfm_3_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_3 <= 1'b0;
    end
    else if ( NMPRun_wen & while_stage_0_4 & (~ while_while_nor_itm_2) ) begin
      while_while_and_itm_3 <= while_while_and_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_2 <= 16'b0000000000000000;
    end
    else if ( NMP_PrepareWriteReq_and_74_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_2 <= NMP_PrepareWriteReq_asn_2_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_2 <= 8'b00000000;
    end
    else if ( NMP_PrepareWriteReq_and_75_enex5 ) begin
      NMP_PrepareWriteReq_asn_1_itm_2 <= NMP_PrepareWriteReq_asn_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_3 <= 2'b00;
    end
    else if ( NMP_PrepareWriteReq_and_53_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_3 <= NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_3 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_3 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_3 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_3_rsp_0 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_3_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_90_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_3 <= rva_out_reg_data_0_sva_dfm_3_2;
      rva_out_reg_data_10_8_sva_dfm_3_3 <= rva_out_reg_data_10_8_sva_dfm_3_2;
      rva_out_reg_data_34_32_sva_dfm_3_3 <= rva_out_reg_data_34_32_sva_dfm_3_2;
      rva_out_reg_data_98_96_sva_dfm_3_3_rsp_0 <= rva_out_reg_data_98_96_sva_dfm_3_2_2;
      rva_out_reg_data_98_96_sva_dfm_3_3_rsp_1 <= rva_out_reg_data_98_96_sva_dfm_3_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_130_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_3 <= rva_out_reg_data_79_64_sva_dfm_3_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_131_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_3 <= rva_out_reg_data_55_48_sva_dfm_3_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_2 <= 1'b0;
    end
    else if ( NMPRun_wen & (~ while_while_nor_itm_1) & while_stage_0_3 ) begin
      while_while_and_itm_2 <= while_while_and_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_1 <= 16'b0000000000000000;
    end
    else if ( NMP_PrepareWriteReq_and_76_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_1 <= nmp_config_timestep_counter_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_1 <= 8'b00000000;
    end
    else if ( NMP_PrepareWriteReq_and_77_enex5 ) begin
      NMP_PrepareWriteReq_asn_1_itm_1 <= nmp_config_vector_counter_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_2 <= 2'b00;
    end
    else if ( NMP_PrepareWriteReq_and_56_cse ) begin
      NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_2 <= reg_nmp_config_adpbias_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3_2 <= 1'b0;
      rva_out_reg_data_10_8_sva_dfm_3_2 <= 3'b000;
      rva_out_reg_data_34_32_sva_dfm_3_2 <= 3'b000;
      rva_out_reg_data_98_96_sva_dfm_3_2_2 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_2_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_96_cse ) begin
      rva_out_reg_data_0_sva_dfm_3_2 <= rva_out_reg_data_0_sva;
      rva_out_reg_data_10_8_sva_dfm_3_2 <= rva_out_reg_data_10_8_sva;
      rva_out_reg_data_34_32_sva_dfm_3_2 <= rva_out_reg_data_34_32_sva;
      rva_out_reg_data_98_96_sva_dfm_3_2_2 <= rva_out_reg_data_98_96_sva_dfm_3_1_2;
      rva_out_reg_data_98_96_sva_dfm_3_2_1_0 <= rva_out_reg_data_98_96_sva_dfm_3_1_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_3_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_132_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_3_2 <= rva_out_reg_data_79_64_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_3_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_133_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_3_2 <= rva_out_reg_data_55_48_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_while_and_itm_1 <= 1'b0;
    end
    else if ( NMPRun_wen & or_503_cse & reg_rva_in_PopNB_mioi_iswt0_cse ) begin
      while_while_and_itm_1 <= NMP_RunFSM_switch_lp_equal_tmp_13 & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva <= 1'b0;
    end
    else if ( NMPRun_wen & (~((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b1100)))
        | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | nand_7_cse)) ) begin
      rva_out_reg_data_0_sva <= nmp_config_is_valid_sva & (~ nmp_config_ConfigRead_unequal_tmp_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_10_8_sva <= 3'b000;
      rva_out_reg_data_79_64_sva <= 16'b0000000000000000;
      rva_out_reg_data_34_32_sva <= 3'b000;
      rva_out_reg_data_55_48_sva <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_1_cse ) begin
      rva_out_reg_data_10_8_sva <= MUX_v_3_2_2(3'b000, nmp_config_mode_sva, nmp_config_ConfigRead_not_12_nl);
      rva_out_reg_data_79_64_sva <= MUX_v_16_2_2(16'b0000000000000000, nmp_config_num_timestep_1_sva,
          nmp_config_ConfigRead_not_10_nl);
      rva_out_reg_data_34_32_sva <= MUX_v_3_2_2(3'b000, nmp_config_memory_index_1_sva,
          nmp_config_ConfigRead_not_9_nl);
      rva_out_reg_data_55_48_sva <= MUX_v_8_2_2(8'b00000000, nmp_config_num_vector_1_sva,
          nmp_config_ConfigRead_not_6_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_1_itm_1_12_9
          <= 4'b0000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_1_itm_1_12_9
          <= MUX_v_4_2_2(ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_12_9,
          (ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_itm_35_11_1[24:21]),
          ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4[0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_1_itm_1_8_0
          <= 9'b000000000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_3_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_1_itm_1_8_0
          <= MUX_v_9_2_2(ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_8_0,
          (ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_itm_35_11_1[20:12]),
          ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4[0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_2_itm_1_10_7
          <= 4'b0000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_4_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_2_itm_1_10_7
          <= MUX_v_4_2_2(ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_7,
          (ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_itm_35_11_1[11:8]),
          ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4[0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_2_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_5_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_mux_2_itm_1_6_0
          <= MUX_v_7_2_2(ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_6_0,
          (ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_temp_mul_itm_35_11_1[7:1]),
          ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4[0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_12_9
          <= 4'b0000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_12_9
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_acc_itm[12:9];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_8_0
          <= 9'b000000000;
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_6_0
          <= 7'b0000000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_8_0
          <= MUX_v_9_2_2((ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_acc_itm[8:0]),
          (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z[42:34]),
          NMP_RunFSM_switch_lp_conc_itm_7_1);
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_6_0
          <= MUX1HOT_v_7_5_2((ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1[6:0]),
          7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, {(~ NMP_RunFSM_switch_lp_conc_itm_7_1)
          , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_nl
          , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_1_nl
          , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_2_nl
          , ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_3_nl});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_7
          <= 4'b0000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_7
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1[10:7];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_2
          <= 1'b0;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_1_0
          <= 2'b00;
    end
    else if ( ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_29_ssc
        ) begin
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_2
          <= (ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_nl
          & (~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_cse)) |
          ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_1_cse | ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_2_cse
          | ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_3_cse;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_1_0
          <= MUX_v_2_2_2(ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_8_nl,
          2'b11, ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_14_itm_1_2
          <= 1'b0;
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_14_itm_1_1_0
          <= 2'b00;
      NMP_PrepareWriteReq_asn_2_itm_7_6_0 <= 7'b0000000;
      NMP_PrepareWriteReq_asn_1_itm_7_7 <= 1'b0;
      NMP_PrepareWriteReq_asn_1_itm_7_6 <= 1'b0;
      NMP_PrepareWriteReq_asn_1_itm_7_5_0 <= 6'b000000;
    end
    else if ( ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_36_ssc
        ) begin
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_14_itm_1_2
          <= (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[33:32]!=2'b00);
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_14_itm_1_1_0
          <= MUX_v_2_2_2(ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_4_nl,
          2'b11, ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_7_cse);
      NMP_PrepareWriteReq_asn_2_itm_7_6_0 <= MUX1HOT_v_7_5_2((NMP_PrepareWriteReq_asn_2_itm_6[6:0]),
          7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, {(~ NMP_RunFSM_switch_lp_conc_itm_7_2)
          , NMP_PrepareWriteReq_and_nl , NMP_PrepareWriteReq_and_1_nl , NMP_PrepareWriteReq_and_2_nl
          , NMP_PrepareWriteReq_and_3_nl});
      NMP_PrepareWriteReq_asn_1_itm_7_7 <= NMP_PrepareWriteReq_asn_1_itm_6_7_6[1];
      NMP_PrepareWriteReq_asn_1_itm_7_6 <= ((NMP_PrepareWriteReq_asn_1_itm_6_7_6[0])
          & (~(NMP_PrepareWriteReq_and_6_ssc | NMP_PrepareWriteReq_and_7_ssc))) |
          NMP_PrepareWriteReq_and_4_ssc | NMP_PrepareWriteReq_and_5_ssc;
      NMP_PrepareWriteReq_asn_1_itm_7_5_0 <= MUX_v_6_2_2(6'b000000, NMP_PrepareWriteReq_NMP_PrepareWriteReq_mux1h_1_nl,
          NMP_PrepareWriteReq_not_6_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_11_8
          <= 4'b0000;
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_7_6
          <= 2'b00;
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_5_0
          <= 6'b000000;
      NMP_PrepareReadReq_asn_2_itm_5_9_0 <= 10'b0000000000;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc
        ) begin
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_11_8
          <= operator_40_0_false_AC_TRN_AC_WRAP_lshift_itm[36:33];
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_7_6
          <= MUX_v_2_2_2(NMP_PrepareReadReq_asn_1_itm_4_7_6, (operator_40_0_false_AC_TRN_AC_WRAP_lshift_itm[32:31]),
          NMP_RunFSM_switch_lp_conc_itm_5_2);
      ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_5_0
          <= MUX_v_6_2_2(NMP_PrepareReadReq_asn_1_itm_4_5_0, (operator_40_0_false_AC_TRN_AC_WRAP_lshift_itm[30:25]),
          NMP_RunFSM_switch_lp_conc_itm_5_2);
      NMP_PrepareReadReq_asn_2_itm_5_9_0 <= MUX1HOT_v_10_5_2((NMP_PrepareReadReq_asn_2_itm_4[9:0]),
          10'b0110101001, 10'b1001010100, 10'b1011101110, 10'b1101111100, {(~ NMP_RunFSM_switch_lp_conc_itm_5_2)
          , NMP_PrepareWriteReq_and_8_cse , NMP_PrepareWriteReq_and_9_cse , NMP_PrepareWriteReq_and_10_cse
          , NMP_PrepareWriteReq_and_11_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_13_rsp_1 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_63_enex5 ) begin
      NMP_PrepareReadReq_asn_1_itm_13_rsp_1 <= NMP_PrepareReadReq_asn_1_itm_12_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_2_36_27 <= 10'b0000000000;
    end
    else if ( NMP_ComputeRMSSqrtRecip_variance_and_enex5 ) begin
      NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_2_36_27 <= NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_36_27;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_2_26_0 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSSqrtRecip_variance_and_2_enex5 ) begin
      NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_2_26_0 <= NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_26_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_36_27 <= 10'b0000000000;
      NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_26_0 <= 27'b000000000000000000000000000;
    end
    else if ( NMP_ComputeRMSSqrtRecip_variance_and_1_ssc ) begin
      NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_36_27 <= NMP_ComputeRMSSqrtRecip_variance_acc_itm[36:27];
      NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_26_0 <= MUX_v_27_2_2((NMP_ComputeRMSSqrtRecip_variance_acc_itm[26:0]),
          NMP_ComputeSoftmaxExp_for_asn_16_itm_2, NMP_RunFSM_switch_lp_conc_itm_3_0);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_12_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_64_enex5 ) begin
      NMP_PrepareReadReq_asn_1_itm_12_5_0 <= NMP_PrepareReadReq_asn_1_itm_11_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_11_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_65_enex5 ) begin
      NMP_PrepareReadReq_asn_1_itm_11_5_0 <= NMP_PrepareReadReq_asn_1_itm_10_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_9_rsp_0 <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_78_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_9_rsp_0 <= NMP_PrepareWriteReq_asn_2_itm_8_15_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_9_rsp_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareWriteReq_and_79_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_9_rsp_1 <= NMP_PrepareWriteReq_asn_2_itm_8_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_0 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_1 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_7_ssc ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_0 <= out_adp_set_value_ac_float_1_asn_15_itm_8_2;
      out_adp_set_value_ac_float_1_asn_15_itm_9_rsp_1 <= out_adp_set_value_ac_float_1_asn_15_itm_8_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_9_rsp_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareReadReq_and_66_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_9_rsp_1 <= NMP_PrepareReadReq_asn_2_itm_8_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_8_15_7 <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_80_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_8_15_7 <= NMP_PrepareWriteReq_asn_2_itm_7_15_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_8_6_0 <= 7'b0000000;
    end
    else if ( NMP_PrepareWriteReq_and_81_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_8_6_0 <= NMP_PrepareWriteReq_asn_2_itm_7_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_8_2 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_8_1_0 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_8_ssc ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_8_2 <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_2;
      out_adp_set_value_ac_float_1_asn_15_itm_8_1_0 <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_10_itm_1_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_8_6_0 <= 7'b0000000;
    end
    else if ( NMP_PrepareReadReq_and_67_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_8_6_0 <= NMP_PrepareReadReq_asn_2_itm_7_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_7_15_7 <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_82_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_7_15_7 <= NMP_PrepareWriteReq_asn_2_itm_6[15:7];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_7_ftd <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_68_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_7_ftd <= NMP_PrepareReadReq_asn_2_itm_6_15_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_7_ftd_1 <= 3'b000;
      NMP_PrepareReadReq_asn_2_itm_7_6_0 <= 7'b0000000;
      NMP_PrepareReadReq_asn_1_itm_7_7 <= 1'b0;
      NMP_PrepareReadReq_asn_1_itm_7_6 <= 1'b0;
      NMP_PrepareReadReq_asn_1_itm_7_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_40_ssc ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_7_ftd_1 <= NMP_PrepareReadReq_asn_2_itm_6_9_0[9:7];
      NMP_PrepareReadReq_asn_2_itm_7_6_0 <= MUX1HOT_v_7_5_2((NMP_PrepareReadReq_asn_2_itm_6_9_0[6:0]),
          7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, {(~ NMP_RunFSM_switch_lp_conc_itm_7_2)
          , NMP_PrepareReadReq_and_2_nl , NMP_PrepareReadReq_and_3_nl , NMP_PrepareReadReq_and_4_nl
          , NMP_PrepareReadReq_and_5_nl});
      NMP_PrepareReadReq_asn_1_itm_7_7 <= NMP_PrepareReadReq_asn_1_itm_6_rsp_0[1];
      NMP_PrepareReadReq_asn_1_itm_7_6 <= ((NMP_PrepareReadReq_asn_1_itm_6_rsp_0[0])
          & (~(ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_5_cse
          | ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_6_cse)))
          | ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_7_cse
          | NMP_PrepareReadReq_and_7_ssc;
      NMP_PrepareReadReq_asn_1_itm_7_5_0 <= MUX_v_6_2_2(6'b000000, NMP_PrepareReadReq_NMP_PrepareReadReq_mux1h_1_nl,
          NMP_PrepareReadReq_not_6_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_6_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_83_enex5 ) begin
      NMP_PrepareWriteReq_asn_1_itm_6_5_0 <= NMP_PrepareWriteReq_asn_1_itm_5_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_6_15_10 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_69_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_6_15_10 <= NMP_PrepareReadReq_asn_2_itm_5_15_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_6_9_0 <= 10'b0000000000;
    end
    else if ( NMP_PrepareReadReq_and_70_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_6_9_0 <= NMP_PrepareReadReq_asn_2_itm_5_9_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_6_rsp_1 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_71_enex5 ) begin
      NMP_PrepareReadReq_asn_1_itm_6_rsp_1 <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_5_7_6 <= 2'b00;
      NMP_PrepareWriteReq_asn_1_itm_5_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_45_ssc ) begin
      NMP_PrepareWriteReq_asn_1_itm_5_7_6 <= NMP_PrepareWriteReq_asn_1_itm_4[7:6];
      NMP_PrepareWriteReq_asn_1_itm_5_5_0 <= MUX1HOT_v_6_5_2((NMP_PrepareWriteReq_asn_1_itm_4[5:0]),
          6'b101011, 6'b011010, 6'b001110, 6'b000100, {(~ NMP_RunFSM_switch_lp_conc_itm_5_2)
          , NMP_PrepareWriteReq_and_8_cse , NMP_PrepareWriteReq_and_9_cse , NMP_PrepareWriteReq_and_10_cse
          , NMP_PrepareWriteReq_and_11_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_5_15_10 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_72_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_5_15_10 <= NMP_PrepareReadReq_asn_2_itm_4[15:10];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_4_7_6 <= 2'b00;
      NMP_PrepareReadReq_asn_1_itm_4_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_48_ssc ) begin
      NMP_PrepareReadReq_asn_1_itm_4_7_6 <= NMP_PrepareReadReq_asn_1_itm_3[7:6];
      NMP_PrepareReadReq_asn_1_itm_4_5_0 <= MUX_v_6_2_2((NMP_PrepareReadReq_asn_1_itm_3[5:0]),
          leading_sign_40_0_out_1, NMP_RunFSM_switch_lp_conc_itm_4_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_3_rsp_0 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_3_rsp_1 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_12_ssc ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_3_rsp_0 <= out_adp_set_value_ac_float_1_asn_15_itm_2_2;
      out_adp_set_value_ac_float_1_asn_15_itm_3_rsp_1 <= out_adp_set_value_ac_float_1_asn_15_itm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_asn_15_itm_3_rsp_0 <= 1'b0;
      out_adp_set_value_ac_float_asn_15_itm_3_rsp_1 <= 2'b00;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_143_cse ) begin
      out_adp_set_value_ac_float_asn_15_itm_3_rsp_0 <= out_adp_set_value_ac_float_1_asn_15_itm_2_2;
      out_adp_set_value_ac_float_asn_15_itm_3_rsp_1 <= out_adp_set_value_ac_float_1_asn_15_itm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_2_2 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_2_1_0 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_13_ssc ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_2_2 <= out_adp_set_value_ac_float_1_asn_15_itm_1_2;
      out_adp_set_value_ac_float_1_asn_15_itm_2_1_0 <= out_adp_set_value_ac_float_1_asn_15_itm_1_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_1_2 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_1_1_0 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_14_ssc ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_1_2 <= reg_nmp_config_adpbias_1_ftd;
      out_adp_set_value_ac_float_1_asn_15_itm_1_1_0 <= reg_nmp_config_adpbias_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_98_96_sva_dfm_3_1_2 <= 1'b0;
      rva_out_reg_data_98_96_sva_dfm_3_1_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_5_ssc ) begin
      rva_out_reg_data_98_96_sva_dfm_3_1_2 <= MUX_s_1_2_2(nmp_config_adpbias_1_sva_dfm_3_1_2,
          nmp_config_ConfigRead_nmp_config_ConfigRead_and_7_nl, while_and_142_rgt);
      rva_out_reg_data_98_96_sva_dfm_3_1_1_0 <= MUX_v_2_2_2(nmp_config_adpbias_1_sva_dfm_3_1_1_0,
          nmp_config_ConfigRead_nmp_config_ConfigRead_and_12_nl, while_and_142_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_16_rsp_1 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_73_enex5 ) begin
      NMP_PrepareReadReq_asn_1_itm_16_rsp_1 <= NMP_PrepareReadReq_asn_1_itm_15_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_15_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_74_enex5 ) begin
      NMP_PrepareReadReq_asn_1_itm_15_5_0 <= reg_NMP_PrepareReadReq_asn_1_itm_14_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_12_rsp_0 <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_84_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_12_rsp_0 <= NMP_PrepareWriteReq_asn_2_itm_11_15_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_12_rsp_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareWriteReq_and_85_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_12_rsp_1 <= NMP_PrepareWriteReq_asn_2_itm_11_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_12_1_ftd_1 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_86_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_12_1_ftd_1 <= NMP_PrepareWriteReq_asn_1_itm_11_6_0_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_12_rsp_0 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_12_rsp_1 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_4_ssc ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_12_rsp_0 <= out_adp_set_value_ac_float_1_asn_15_itm_11_2;
      out_adp_set_value_ac_float_1_asn_15_itm_12_rsp_1 <= out_adp_set_value_ac_float_1_asn_15_itm_11_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_asn_15_itm_12_rsp_0 <= 1'b0;
      out_adp_set_value_ac_float_asn_15_itm_12_rsp_1 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_and_4_ssc ) begin
      out_adp_set_value_ac_float_asn_15_itm_12_rsp_0 <= out_adp_set_value_ac_float_asn_15_itm_11_2;
      out_adp_set_value_ac_float_asn_15_itm_12_rsp_1 <= out_adp_set_value_ac_float_asn_15_itm_11_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_12_ftd <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_75_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_12_ftd <= NMP_PrepareReadReq_asn_2_itm_11_15_7_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_12_rsp_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareReadReq_and_76_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_12_rsp_1 <= NMP_PrepareReadReq_asn_2_itm_11_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_11_15_7 <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_87_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_11_15_7 <= reg_NMP_PrepareWriteReq_asn_2_itm_10_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_11_6_0 <= 7'b0000000;
    end
    else if ( NMP_PrepareWriteReq_and_88_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_11_6_0 <= reg_NMP_PrepareWriteReq_asn_2_itm_10_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_11_2 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_11_1_0 <= 2'b00;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_cse ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_11_2 <= reg_out_adp_set_value_ac_float_1_asn_15_itm_10_ftd;
      out_adp_set_value_ac_float_1_asn_15_itm_11_1_0 <= reg_out_adp_set_value_ac_float_1_asn_15_itm_10_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_asn_15_itm_11_2 <= 1'b0;
      out_adp_set_value_ac_float_asn_15_itm_11_1_0 <= 2'b00;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_cse ) begin
      out_adp_set_value_ac_float_asn_15_itm_11_2 <= reg_out_adp_set_value_ac_float_asn_15_itm_10_ftd;
      out_adp_set_value_ac_float_asn_15_itm_11_1_0 <= reg_out_adp_set_value_ac_float_asn_15_itm_10_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_11_6_0 <= 7'b0000000;
    end
    else if ( NMP_PrepareReadReq_and_77_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_11_6_0 <= reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_6_rsp_0 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_6_rsp_1 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_9_ssc ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_6_rsp_0 <= out_adp_set_value_ac_float_1_asn_15_itm_5_2;
      out_adp_set_value_ac_float_1_asn_15_itm_6_rsp_1 <= out_adp_set_value_ac_float_1_asn_15_itm_5_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_asn_15_itm_6_rsp_0 <= 1'b0;
      out_adp_set_value_ac_float_asn_15_itm_6_rsp_1 <= 2'b00;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_96_cse ) begin
      out_adp_set_value_ac_float_asn_15_itm_6_rsp_0 <= out_adp_set_value_ac_float_asn_15_itm_5_2;
      out_adp_set_value_ac_float_asn_15_itm_6_rsp_1 <= out_adp_set_value_ac_float_asn_15_itm_5_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_5_2 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_5_1_0 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_10_ssc ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_5_2 <= reg_out_adp_set_value_ac_float_1_asn_15_itm_4_ftd;
      out_adp_set_value_ac_float_1_asn_15_itm_5_1_0 <= reg_out_adp_set_value_ac_float_1_asn_15_itm_4_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_asn_15_itm_5_2 <= 1'b0;
      out_adp_set_value_ac_float_asn_15_itm_5_1_0 <= 2'b00;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_112_cse ) begin
      out_adp_set_value_ac_float_asn_15_itm_5_2 <= reg_out_adp_set_value_ac_float_asn_15_itm_4_ftd;
      out_adp_set_value_ac_float_asn_15_itm_5_1_0 <= reg_out_adp_set_value_ac_float_asn_15_itm_4_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_9_rsp_1_rsp_1 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_89_enex5 ) begin
      NMP_PrepareWriteReq_asn_1_itm_9_rsp_1_rsp_1 <= NMP_PrepareWriteReq_asn_1_itm_8_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_9_rsp_0_rsp_0 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_78_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_9_rsp_0_rsp_0 <= NMP_PrepareReadReq_asn_2_itm_8_15_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_9_rsp_1_rsp_1 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_79_enex5 ) begin
      NMP_PrepareReadReq_asn_1_itm_9_rsp_1_rsp_1 <= NMP_PrepareReadReq_asn_1_itm_8_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_8_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_90_enex5 ) begin
      NMP_PrepareWriteReq_asn_1_itm_8_5_0 <= NMP_PrepareWriteReq_asn_1_itm_7_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_8_15_10 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_80_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_8_15_10 <= reg_NMP_PrepareReadReq_asn_2_itm_7_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_1_itm_8_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_81_enex5 ) begin
      NMP_PrepareReadReq_asn_1_itm_8_5_0 <= NMP_PrepareReadReq_asn_1_itm_7_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_15_rsp_0 <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_91_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_15_rsp_0 <= NMP_PrepareWriteReq_asn_2_itm_14_15_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_15_rsp_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareWriteReq_and_92_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_15_rsp_1 <= NMP_PrepareWriteReq_asn_2_itm_14_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_15_1_ftd_1 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_93_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_15_1_ftd_1 <= NMP_PrepareWriteReq_asn_1_itm_14_6_0_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_15_ftd <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_82_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_15_ftd <= NMP_PrepareReadReq_asn_2_itm_14_15_7_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_15_rsp_1 <= 7'b0000000;
    end
    else if ( NMP_PrepareReadReq_and_83_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_15_rsp_1 <= NMP_PrepareReadReq_asn_2_itm_14_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_14_15_7 <= 9'b000000000;
    end
    else if ( NMP_PrepareWriteReq_and_94_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_14_15_7 <= reg_NMP_PrepareWriteReq_asn_2_itm_13_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_2_itm_14_6_0 <= 7'b0000000;
    end
    else if ( NMP_PrepareWriteReq_and_95_enex5 ) begin
      NMP_PrepareWriteReq_asn_2_itm_14_6_0 <= reg_NMP_PrepareWriteReq_asn_2_itm_13_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_14_2 <= 1'b0;
      out_adp_set_value_ac_float_1_asn_15_itm_14_1_0 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_1_and_2_ssc ) begin
      out_adp_set_value_ac_float_1_asn_15_itm_14_2 <= reg_out_adp_set_value_ac_float_1_asn_15_itm_13_ftd;
      out_adp_set_value_ac_float_1_asn_15_itm_14_1_0 <= reg_out_adp_set_value_ac_float_1_asn_15_itm_13_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      out_adp_set_value_ac_float_asn_15_itm_14_2 <= 1'b0;
      out_adp_set_value_ac_float_asn_15_itm_14_1_0 <= 2'b00;
    end
    else if ( out_adp_set_value_ac_float_and_2_ssc ) begin
      out_adp_set_value_ac_float_asn_15_itm_14_2 <= reg_out_adp_set_value_ac_float_asn_15_itm_13_ftd;
      out_adp_set_value_ac_float_asn_15_itm_14_1_0 <= reg_out_adp_set_value_ac_float_asn_15_itm_13_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_14_6_0 <= 7'b0000000;
    end
    else if ( NMP_PrepareReadReq_and_84_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_14_6_0 <= reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_11_6_0_rsp_1 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_96_enex5 ) begin
      NMP_PrepareWriteReq_asn_1_itm_11_6_0_rsp_1 <= reg_NMP_PrepareWriteReq_asn_1_itm_10_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_11_15_7_rsp_0 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_85_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_11_15_7_rsp_0 <= reg_NMP_PrepareReadReq_asn_2_itm_10_ftd_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd_1_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_97_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd_1_5_0 <= reg_NMP_PrepareWriteReq_asn_1_itm_12_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_8_3 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_86_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_8_3 <= reg_NMP_PrepareReadReq_asn_2_itm_12_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareWriteReq_asn_1_itm_14_6_0_rsp_1 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_98_enex5 ) begin
      NMP_PrepareWriteReq_asn_1_itm_14_6_0_rsp_1 <= reg_NMP_PrepareWriteReq_asn_1_itm_13_ftd_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      NMP_PrepareReadReq_asn_2_itm_14_15_7_rsp_0 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_87_enex5 ) begin
      NMP_PrepareReadReq_asn_2_itm_14_15_7_rsp_0 <= reg_NMP_PrepareReadReq_asn_2_itm_13_ftd_8_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_8_3 <= 6'b000000;
    end
    else if ( NMP_PrepareReadReq_and_88_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_16_ftd_8_3 <= reg_NMP_PrepareReadReq_asn_2_itm_15_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd_1_5_0 <= 6'b000000;
    end
    else if ( NMP_PrepareWriteReq_and_99_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_16_ftd_1_5_0 <= reg_NMP_PrepareWriteReq_asn_1_itm_15_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_15_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_16_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_15_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_1_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_15_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_16_enex5
        ) begin
      reg_out_float_round_32_if_m_1_1_sva_1_6_enexo <= out_float_round_32_if_m_1_and_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_16_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_16_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_1_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_31_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_16_enex5
        ) begin
      reg_out_float_round_32_if_m_1_1_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_31_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_15_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_16_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_15_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_1_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_31_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_16_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_1_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_31_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_1_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_15_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_16_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_1_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_16_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_16_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_17_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_14_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_17_enex5
        ) begin
      reg_out_float_round_32_if_m_1_17_sva_1_6_enexo <= out_float_round_32_if_m_1_and_14_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_17_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_30_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_17_enex5
        ) begin
      reg_out_float_round_32_if_m_1_17_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_30_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_17_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_15_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_17_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_15_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_17_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_14_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_17_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_17_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_14_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_17_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_15_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_14_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_17_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_14_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_17_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_30_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_17_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_17_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_30_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_13_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_18_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_13_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_18_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_14_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_16_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_29_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_18_enex5
        ) begin
      reg_out_float_round_32_if_m_1_16_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_29_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_16_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_13_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_18_enex5
        ) begin
      reg_out_float_round_32_if_m_1_16_sva_1_6_enexo <= out_float_round_32_if_m_1_and_13_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_18_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_14_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_18_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_14_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_16_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_29_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_18_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_16_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_29_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_16_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_13_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_18_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_16_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_13_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_15_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_12_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_19_enex5
        ) begin
      reg_out_float_round_32_if_m_1_15_sva_1_6_enexo <= out_float_round_32_if_m_1_and_12_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_3 <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_19_enex5
        ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_3 <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_15_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_28_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_19_enex5
        ) begin
      reg_out_float_round_32_if_m_1_15_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_28_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_19_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_13_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_12_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_19_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_12_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_15_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_12_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_19_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_15_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_12_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_19_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_13_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_15_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_28_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_19_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_15_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_28_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_20_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_12_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_14_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_27_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_20_enex5
        ) begin
      reg_out_float_round_32_if_m_1_14_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_27_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_14_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_11_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_20_enex5
        ) begin
      reg_out_float_round_32_if_m_1_14_sva_1_6_enexo <= out_float_round_32_if_m_1_and_11_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_20_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_12_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_20_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_12_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_14_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_27_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_20_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_14_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_27_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_11_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_20_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_11_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_14_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_11_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_20_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_14_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_11_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_13_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_26_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_21_enex5
        ) begin
      reg_out_float_round_32_if_m_1_13_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_26_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_13_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_10_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_21_enex5
        ) begin
      reg_out_float_round_32_if_m_1_13_sva_1_6_enexo <= out_float_round_32_if_m_1_and_10_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_21_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_11_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_21_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_11_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_10_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_21_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_10_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_13_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_10_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_21_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_13_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_10_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_13_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_26_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_21_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_13_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_26_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_21_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_11_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_22_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_10_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_22_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_10_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_12_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_25_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_22_enex5
        ) begin
      reg_out_float_round_32_if_m_1_12_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_25_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_12_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_9_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_22_enex5
        ) begin
      reg_out_float_round_32_if_m_1_12_sva_1_6_enexo <= out_float_round_32_if_m_1_and_9_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_22_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_10_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_22_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_10_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_12_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_25_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_22_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_12_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_25_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_12_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_9_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_22_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_12_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_9_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_11_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_24_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_23_enex5
        ) begin
      reg_out_float_round_32_if_m_1_11_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_24_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_23_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_9_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_7 <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_23_enex5
        ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_7 <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_11_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_8_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_23_enex5
        ) begin
      reg_out_float_round_32_if_m_1_11_sva_1_6_enexo <= out_float_round_32_if_m_1_and_8_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_8_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_23_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_8_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_23_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_9_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_11_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_8_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_23_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_11_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_8_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_11_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_24_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_23_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_11_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_24_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_10_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_7_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_24_enex5
        ) begin
      reg_out_float_round_32_if_m_1_10_sva_1_6_enexo <= out_float_round_32_if_m_1_and_7_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_24_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_8_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_24_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_8_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_10_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_23_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_24_enex5
        ) begin
      reg_out_float_round_32_if_m_1_10_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_23_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_24_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_8_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_24_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_8_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_10_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_23_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_24_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_10_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_23_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_10_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_7_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_24_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_10_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_7_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_9_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_22_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_25_enex5
        ) begin
      reg_out_float_round_32_if_m_1_9_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_22_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_6_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_25_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_6_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_9_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_6_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_25_enex5
        ) begin
      reg_out_float_round_32_if_m_1_9_sva_1_6_enexo <= out_float_round_32_if_m_1_and_6_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_25_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_7_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_6_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_25_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_6_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_9_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_22_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_25_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_9_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_22_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_25_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_7_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_9_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_6_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_25_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_9_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_6_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_26_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_6_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_8_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_21_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_26_enex5
        ) begin
      reg_out_float_round_32_if_m_1_8_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_21_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_8_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_5_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_26_enex5
        ) begin
      reg_out_float_round_32_if_m_1_8_sva_1_6_enexo <= out_float_round_32_if_m_1_and_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_26_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_6_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_26_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_6_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_8_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_21_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_26_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_8_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_21_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_8_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_5_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_26_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_8_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_26_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_6_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_27_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_5_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_27_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_eq_in_ac_float_compare_32_32_1_AC_TRN_eq_nor_5_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_7_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_20_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_27_enex5
        ) begin
      reg_out_float_round_32_if_m_1_7_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_20_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_7_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_4_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_27_enex5
        ) begin
      reg_out_float_round_32_if_m_1_7_sva_1_6_enexo <= out_float_round_32_if_m_1_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_7_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_4_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_27_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_7_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_4_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_27_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_and_4_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_27_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_5_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_7_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_20_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_27_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_7_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_20_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_6_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_19_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_28_enex5
        ) begin
      reg_out_float_round_32_if_m_1_6_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_19_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_3_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_28_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_3_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_6_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_3_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_28_enex5
        ) begin
      reg_out_float_round_32_if_m_1_6_sva_1_6_enexo <= out_float_round_32_if_m_1_and_3_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_28_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_4_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_28_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_4_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_6_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_19_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_28_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_6_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_19_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_6_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_3_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_28_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_6_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_3_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_28_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_4_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_5_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_2_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_29_enex5
        ) begin
      reg_out_float_round_32_if_m_1_5_sva_1_6_enexo <= out_float_round_32_if_m_1_and_2_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_2_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_29_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_2_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_5_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_18_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_29_enex5
        ) begin
      reg_out_float_round_32_if_m_1_5_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_18_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_29_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_3_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_29_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_3_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_5_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_18_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_29_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_5_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_18_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_29_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_3_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_5_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_2_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_29_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_5_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_2_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_4_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_1_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_30_enex5
        ) begin
      reg_out_float_round_32_if_m_1_4_sva_1_6_enexo <= out_float_round_32_if_m_1_and_1_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_14 <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_30_enex5
        ) begin
      reg_out_adp_set_value_ac_float_asn_15_itm_16_enexo_14 <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_4_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_17_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_30_enex5
        ) begin
      reg_out_float_round_32_if_m_1_4_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_17_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_30_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_2_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_30_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_2_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_4_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_1_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_30_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_4_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_1_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_30_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_2_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_4_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_17_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_30_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_4_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_17_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_3_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_31_enex5
        ) begin
      reg_out_float_round_32_if_m_1_3_sva_1_6_enexo <= out_float_round_32_if_m_1_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_if_m_1_3_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_if_m_1_and_16_tmp | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_31_enex5
        ) begin
      reg_out_float_round_32_if_m_1_3_sva_1_3_0_enexo <= out_float_round_32_if_m_1_and_16_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_31_enex5
        ) begin
      reg_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_and_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_and_cse | NMP_ConvertOutputToAdpfloat_for_out_adp_man_and_31_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_for_1_operator_6_2_true_AC_TRN_AC_WRAP_operator_6_2_true_AC_TRN_AC_WRAP_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= 1'b1;
    end
    else if ( operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_31_enex5
        ) begin
      reg_NMP_ConvertOutputToAdpfloat_1_for_1_operator_6_2_true_AC_TRN_AC_WRAP_1_operator_6_2_true_AC_TRN_AC_WRAP_1_and_svs_enexo
          <= operator_6_2_true_AC_TRN_AC_WRAP_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_3_sva_1_3_0_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_16_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_31_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_3_sva_1_3_0_enexo <= out_float_round_32_1_if_m_1_and_16_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1_enexo
          <= 1'b1;
    end
    else if ( in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_31_enex5
        ) begin
      reg_in_ac_float_compare_32_32_1_AC_TRN_1_eq_in_ac_float_compare_32_32_1_AC_TRN_1_eq_nor_itm_1_enexo
          <= in_ac_float_compare_32_32_1_AC_TRN_1_eq_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_out_float_round_32_1_if_m_1_3_sva_1_6_enexo <= 1'b1;
    end
    else if ( out_float_round_32_1_if_m_1_and_tmp | NMP_ConvertOutputToAdpfloat_1_for_out_adp_man_and_31_enex5
        ) begin
      reg_out_float_round_32_1_if_m_1_3_sva_1_6_enexo <= out_float_round_32_1_if_m_1_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_15_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_83_enex5 | NMP_PrepareReadReq_and_55_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_15_1_enexo <= NMP_PrepareReadReq_and_83_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_15_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_91_enex5 | NMP_PrepareWriteReq_and_61_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_15_enexo <= NMP_PrepareWriteReq_and_91_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_15_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_92_enex5 | NMP_PrepareWriteReq_and_62_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_15_1_enexo <= NMP_PrepareWriteReq_and_92_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_16_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_104_enex5 | rva_out_reg_data_and_102_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_16_enexo <= rva_out_reg_data_and_104_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_16_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_105_enex5 | rva_out_reg_data_and_103_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_16_enexo <= rva_out_reg_data_and_105_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_6_enex5
        | ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5
        ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_enexo
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_6_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_3_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_enex5
        | ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_3_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_1_cse
        | ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5
        ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_2_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_4_enex5
        | ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_3_enex5 )
        begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_itm_2_enexo
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_4_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_2_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_2_enex5
        | ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_1_enex5
        ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_itm_2_enexo
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_2_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_1_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_2_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_1_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_161_enex5 | NMP_ComputeRMSNormalize_for_and_145_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_161_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_162_enex5 | NMP_ComputeRMSNormalize_for_and_146_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_162_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_163_enex5 | NMP_ComputeRMSNormalize_for_and_147_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_163_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_164_enex5 | NMP_ComputeRMSNormalize_for_and_148_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_164_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_165_enex5 | NMP_ComputeRMSNormalize_for_and_149_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_165_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_166_enex5 | NMP_ComputeRMSNormalize_for_and_150_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_166_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_167_enex5 | NMP_ComputeRMSNormalize_for_and_151_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_167_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_168_enex5 | NMP_ComputeRMSNormalize_for_and_152_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_168_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_169_enex5 | NMP_ComputeRMSNormalize_for_and_153_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_169_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_170_enex5 | NMP_ComputeRMSNormalize_for_and_154_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_170_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_171_enex5 | NMP_ComputeRMSNormalize_for_and_155_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_171_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_172_enex5 | NMP_ComputeRMSNormalize_for_and_156_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_172_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_173_enex5 | NMP_ComputeRMSNormalize_for_and_157_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_173_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_10_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_174_enex5 | NMP_ComputeRMSNormalize_for_and_158_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_10_enexo <= NMP_ComputeRMSNormalize_for_and_174_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_10_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_175_enex5 | NMP_ComputeRMSNormalize_for_and_159_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_10_enexo <= NMP_ComputeRMSNormalize_for_and_175_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_10_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_176_enex5 | NMP_ComputeRMSNormalize_for_and_160_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_10_enexo <= NMP_ComputeRMSNormalize_for_and_176_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_sum_exp_39_4_sva_st_3_enexo <= 1'b1;
    end
    else if ( sum_exp_and_1_enex5 | sum_exp_and_enex5 ) begin
      reg_sum_exp_39_4_sva_st_3_enexo <= sum_exp_and_1_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_96_enex5 | NMP_ComputeSoftmaxNormalize_for_and_80_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_96_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_97_enex5 | NMP_ComputeSoftmaxNormalize_for_and_81_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_97_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_98_enex5 | NMP_ComputeSoftmaxNormalize_for_and_82_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_98_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_99_enex5 | NMP_ComputeSoftmaxNormalize_for_and_83_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_99_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_100_enex5 | NMP_ComputeSoftmaxNormalize_for_and_84_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_100_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_101_enex5 | NMP_ComputeSoftmaxNormalize_for_and_85_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_101_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_102_enex5 | NMP_ComputeSoftmaxNormalize_for_and_86_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_102_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_103_enex5 | NMP_ComputeSoftmaxNormalize_for_and_87_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_103_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_104_enex5 | NMP_ComputeSoftmaxNormalize_for_and_88_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_104_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_105_enex5 | NMP_ComputeSoftmaxNormalize_for_and_89_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_105_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_106_enex5 | NMP_ComputeSoftmaxNormalize_for_and_90_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_106_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_107_enex5 | NMP_ComputeSoftmaxNormalize_for_and_91_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_107_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_108_enex5 | NMP_ComputeSoftmaxNormalize_for_and_92_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_108_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_109_enex5 | NMP_ComputeSoftmaxNormalize_for_and_93_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_109_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_110_enex5 | NMP_ComputeSoftmaxNormalize_for_and_94_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_110_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_111_enex5 | NMP_ComputeSoftmaxNormalize_for_and_95_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_3_enexo <= NMP_ComputeSoftmaxNormalize_for_and_111_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_1_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_2_cse
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_1_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qr_sva_st_1_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_sum_exp_39_4_sva_st_2_enexo <= 1'b1;
    end
    else if ( sum_exp_and_2_enex5 | sum_exp_and_1_enex5 ) begin
      reg_sum_exp_39_4_sva_st_2_enexo <= sum_exp_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_sum_exp_39_4_sva_st_1_enexo <= 1'b1;
    end
    else if ( sum_exp_and_3_enex5 | sum_exp_and_2_enex5 ) begin
      reg_sum_exp_39_4_sva_st_1_enexo <= sum_exp_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp |
        ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_12_enex5 ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_50_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_50_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_50_enex5 ) begin
      reg_max_value_26_0_1_enexo <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_50_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_30_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_66_enex5 | NMP_ComputeSoftmaxExp_for_and_50_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_30_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_50_enex5 ) begin
      reg_while_stage_0_7_enexo <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_50_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_50_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_50_enex5 ) begin
      reg_max_value_26_0_enexo <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_1 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_51_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_1 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_67_enex5 | NMP_ComputeSoftmaxExp_for_and_51_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_1 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_51_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_1 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_1 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_51_enex5 ) begin
      reg_max_value_26_0_1_enexo_1 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_1 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_51_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_1 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_1 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_51_enex5 ) begin
      reg_while_stage_0_7_enexo_1 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_51_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_1 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_1 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_51_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_1 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_1 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_51_enex5 ) begin
      reg_max_value_26_0_enexo_1 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_2 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_52_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_2 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_2 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_52_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_2 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_2 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_52_enex5 ) begin
      reg_max_value_26_0_1_enexo_2 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_2 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_52_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_2 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_2 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_52_enex5 ) begin
      reg_while_stage_0_7_enexo_2 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_2 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_52_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_2 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_2 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_52_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_2 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_2 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_52_enex5 ) begin
      reg_max_value_26_0_enexo_2 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_68_enex5 | NMP_ComputeSoftmaxExp_for_and_52_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_3 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_53_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_3 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_3 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_53_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_3 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_3 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_53_enex5 ) begin
      reg_max_value_26_0_1_enexo_3 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_69_enex5 | NMP_ComputeSoftmaxExp_for_and_53_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_3 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_53_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_3 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_3 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_53_enex5 ) begin
      reg_while_stage_0_7_enexo_3 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_3 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_53_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_3 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_3 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_53_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_3 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_3 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_53_enex5 ) begin
      reg_max_value_26_0_enexo_3 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_4 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_54_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_4 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_70_enex5 | NMP_ComputeSoftmaxExp_for_and_54_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_70_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_4 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_54_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_4 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_4 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_54_enex5 ) begin
      reg_max_value_26_0_1_enexo_4 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_4 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_54_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_4 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_4 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_54_enex5 ) begin
      reg_while_stage_0_7_enexo_4 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_4 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_54_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_4 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_4 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_54_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_4 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_4 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_54_enex5 ) begin
      reg_max_value_26_0_enexo_4 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_5 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_55_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_5 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_5 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_55_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_5 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_5 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_55_enex5 ) begin
      reg_max_value_26_0_1_enexo_5 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_5 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_55_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_5 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_5 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_55_enex5 ) begin
      reg_while_stage_0_7_enexo_5 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_5 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_55_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_5 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_5 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_55_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_5 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_5 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_55_enex5 ) begin
      reg_max_value_26_0_enexo_5 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_21_enex5 | NMP_ComputeSoftmaxExp_for_and_55_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_6 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_56_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_6 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_71_enex5 | NMP_ComputeSoftmaxExp_for_and_56_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_71_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_6 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_56_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_6 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_6 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_56_enex5 ) begin
      reg_max_value_26_0_1_enexo_6 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_6 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_56_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_6 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_6 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_56_enex5 ) begin
      reg_while_stage_0_7_enexo_6 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_6 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_56_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_6 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_6 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_56_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_6 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_6 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_56_enex5 ) begin
      reg_max_value_26_0_enexo_6 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_7 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_57_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_7 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_7 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_57_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_7 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_7 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_57_enex5 ) begin
      reg_max_value_26_0_1_enexo_7 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_72_enex5 | NMP_ComputeSoftmaxExp_for_and_57_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_72_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_7 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_57_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_7 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_7 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_57_enex5 ) begin
      reg_while_stage_0_7_enexo_7 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_7 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_57_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_7 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_7 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_57_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_7 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_7 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_57_enex5 ) begin
      reg_max_value_26_0_enexo_7 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_8 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_58_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_8 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_73_enex5 | NMP_ComputeSoftmaxExp_for_and_58_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_73_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_8 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_58_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_8 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_8 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_58_enex5 ) begin
      reg_max_value_26_0_1_enexo_8 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_8 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_58_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_8 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_8 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_58_enex5 ) begin
      reg_while_stage_0_7_enexo_8 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_8 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_58_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_8 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_8 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_58_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_8 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_8 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_58_enex5 ) begin
      reg_max_value_26_0_enexo_8 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_9 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_59_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_9 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_9 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_59_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_9 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_9 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_59_enex5 ) begin
      reg_max_value_26_0_1_enexo_9 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_9 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_59_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_9 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_9 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_59_enex5 ) begin
      reg_while_stage_0_7_enexo_9 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_9 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_59_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_9 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_9 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_59_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_9 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_9 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_59_enex5 ) begin
      reg_max_value_26_0_enexo_9 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_74_enex5 | NMP_ComputeSoftmaxExp_for_and_59_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_74_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_10 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_60_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_10 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_10 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_60_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_10 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_10 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_60_enex5 ) begin
      reg_max_value_26_0_1_enexo_10 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_10 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_60_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_10 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_10 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_60_enex5 ) begin
      reg_while_stage_0_7_enexo_10 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_75_enex5 | NMP_ComputeSoftmaxExp_for_and_60_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_75_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_10 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_60_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_10 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_10 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_60_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_10 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_10 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_60_enex5 ) begin
      reg_max_value_26_0_enexo_10 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_11 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_61_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_11 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_76_enex5 | NMP_ComputeSoftmaxExp_for_and_61_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_76_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_11 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_61_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_11 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_11 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_61_enex5 ) begin
      reg_max_value_26_0_1_enexo_11 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_11 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_61_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_11 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_11 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_61_enex5 ) begin
      reg_while_stage_0_7_enexo_11 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_11 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_61_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_11 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_11 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_61_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_11 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_11 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_61_enex5 ) begin
      reg_max_value_26_0_enexo_11 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_12 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_62_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_12 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_12 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_62_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_12 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_12 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_62_enex5 ) begin
      reg_max_value_26_0_1_enexo_12 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_12 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_62_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_12 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_12 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_62_enex5 ) begin
      reg_while_stage_0_7_enexo_12 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_12 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_62_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_12 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_12 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_62_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_12 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_12 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_62_enex5 ) begin
      reg_max_value_26_0_enexo_12 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_77_enex5 | NMP_ComputeSoftmaxExp_for_and_62_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_77_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_78_enex5 | NMP_ComputeSoftmaxExp_for_and_63_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_3_enexo <= NMP_ComputeSoftmaxExp_for_and_78_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_13 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_63_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_13 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_13 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_63_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_13 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_13 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_63_enex5 ) begin
      reg_max_value_26_0_1_enexo_13 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_13 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_63_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_13 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_13 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_63_enex5 ) begin
      reg_while_stage_0_7_enexo_13 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_13 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_63_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_13 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_13 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_63_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_13 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_13 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_63_enex5 ) begin
      reg_max_value_26_0_enexo_13 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_14 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_64_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_14 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_14 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_64_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_14 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_14 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_64_enex5 ) begin
      reg_max_value_26_0_1_enexo_14 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_14 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_64_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_14 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_14 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_64_enex5 ) begin
      reg_while_stage_0_7_enexo_14 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_79_enex5 | NMP_ComputeSoftmaxExp_for_and_64_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_3_enexo <= NMP_ComputeSoftmaxExp_for_and_79_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_14 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_64_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_14 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_14 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_64_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_14 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_14 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_64_enex5 ) begin
      reg_max_value_26_0_enexo_14 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_15 <= 1'b1;
    end
    else if ( while_if_and_13_cse | NMP_ComputeSoftmaxExp_for_and_65_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_15 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_15 <= 1'b1;
    end
    else if ( max_value_and_enex5 | NMP_ComputeSoftmaxExp_for_and_65_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_15 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_15 <= 1'b1;
    end
    else if ( and_1085_enex5 | NMP_ComputeSoftmaxExp_for_and_65_enex5 ) begin
      reg_max_value_26_0_1_enexo_15 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_15 <= 1'b1;
    end
    else if ( max_value_and_1_cse | NMP_ComputeSoftmaxExp_for_and_65_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_15 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_stage_0_7_enexo_15 <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_ComputeSoftmaxExp_for_and_65_enex5 ) begin
      reg_while_stage_0_7_enexo_15 <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_15 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | NMP_ComputeSoftmaxExp_for_and_65_enex5
        ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_15 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_15 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeSoftmaxExp_for_and_65_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_15 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_enexo_15 <= 1'b1;
    end
    else if ( while_if_and_12_cse | NMP_ComputeSoftmaxExp_for_and_65_enex5 ) begin
      reg_max_value_26_0_enexo_15 <= while_if_and_12_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_80_enex5 | NMP_ComputeSoftmaxExp_for_and_65_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_itm_3_enexo <= NMP_ComputeSoftmaxExp_for_and_80_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_1_cse
        | ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_5_enex5
        ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_enexo
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo_2
          <= 1'b1;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_1_cse
        | ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_6_enex5
        ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo_2
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_2_cse
        | ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_4_enex5
        ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_slc_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_normalized_fixed_38_26_9_0_enexo
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_2_cse
        | ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_5_enex5
        ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_enexo
          <= ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_and_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_16 <= 1'b1;
    end
    else if ( while_if_and_13_cse | and_1085_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_equal_tmp_5_4_enexo_16 <= while_if_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_16 <= 1'b1;
    end
    else if ( max_value_and_enex5 | and_1085_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_25_0_enexo_16 <= max_value_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_1_enexo_16 <= 1'b1;
    end
    else if ( and_1085_enex5 ) begin
      reg_max_value_26_0_1_enexo_16 <= and_1085_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_16 <= 1'b1;
    end
    else if ( max_value_and_1_cse | and_1085_enex5 ) begin
      reg_max_value_26_0_sva_dfm_13_1_26_enexo_16 <= max_value_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_16 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_and_enex5 | and_1085_enex5 ) begin
      reg_NMP_ComputeSoftmaxMax_for_asn_13_itm_3_enexo_16 <= NMP_ComputeSoftmaxMax_for_and_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_16 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | and_1085_enex5 ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_16 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_30_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_66_enex5 | NMP_RunFSM_switch_lp_and_126_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_30_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_67_enex5 | NMP_ComputeSoftmaxMax_for_and_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_9_1_25_0_enexo <= 1'b1;
    end
    else if ( max_value_and_9_enex5 | max_value_and_enex5 ) begin
      reg_max_value_26_0_sva_dfm_9_1_25_0_enexo <= max_value_and_9_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxMax_for_if_less_5_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxMax_for_if_and_tmp | max_value_and_enex5 ) begin
      reg_NMP_ComputeSoftmaxMax_for_if_less_5_itm_1_enexo <= NMP_ComputeSoftmaxMax_for_if_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_70_enex5 | max_value_and_enex5 ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_70_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_69_enex5 | max_value_and_enex5 ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_9_1_26_enexo <= 1'b1;
    end
    else if ( max_value_and_3_cse | max_value_and_enex5 ) begin
      reg_max_value_26_0_sva_dfm_9_1_26_enexo <= max_value_and_3_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_68_enex5 | max_value_and_enex5 ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_21_enex5 | max_value_and_enex5 ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_342_enex5 | NMP_ComputeSoftmaxExp_for_and_66_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_1_enexo <= NMP_RunFSM_switch_lp_and_342_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_81_enex5 | NMP_ComputeSoftmaxExp_for_and_67_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_81_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_82_enex5 | NMP_ComputeSoftmaxExp_for_and_68_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_82_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_83_enex5 | NMP_ComputeSoftmaxExp_for_and_69_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_83_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_84_enex5 | NMP_ComputeSoftmaxExp_for_and_70_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_84_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_85_enex5 | NMP_ComputeSoftmaxExp_for_and_21_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_85_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_86_enex5 | NMP_ComputeSoftmaxExp_for_and_71_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_86_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_87_enex5 | NMP_ComputeSoftmaxExp_for_and_72_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_87_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_88_enex5 | NMP_ComputeSoftmaxExp_for_and_73_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_88_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_89_enex5 | NMP_ComputeSoftmaxExp_for_and_74_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_89_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_90_enex5 | NMP_ComputeSoftmaxExp_for_and_75_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_90_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_91_enex5 | NMP_ComputeSoftmaxExp_for_and_76_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_91_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_92_enex5 | NMP_ComputeSoftmaxExp_for_and_77_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_92_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_93_enex5 | NMP_ComputeSoftmaxExp_for_and_78_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_93_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_94_enex5 | NMP_ComputeSoftmaxExp_for_and_79_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_94_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_95_enex5 | NMP_ComputeSoftmaxExp_for_and_80_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_itm_2_enexo <= NMP_ComputeSoftmaxExp_for_and_95_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxSum_for_acc_7_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxSum_for_and_cse | sum_exp_and_3_enex5 ) begin
      reg_NMP_ComputeSoftmaxSum_for_acc_7_itm_1_enexo <= NMP_ComputeSoftmaxSum_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_112_enex5 | NMP_ComputeSoftmaxNormalize_for_and_96_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_112_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_113_enex5 | NMP_ComputeSoftmaxNormalize_for_and_97_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_113_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_114_enex5 | NMP_ComputeSoftmaxNormalize_for_and_98_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_114_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_115_enex5 | NMP_ComputeSoftmaxNormalize_for_and_99_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_115_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_116_enex5 | NMP_ComputeSoftmaxNormalize_for_and_100_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_116_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_117_enex5 | NMP_ComputeSoftmaxNormalize_for_and_101_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_117_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_118_enex5 | NMP_ComputeSoftmaxNormalize_for_and_102_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_118_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_119_enex5 | NMP_ComputeSoftmaxNormalize_for_and_103_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_119_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_120_enex5 | NMP_ComputeSoftmaxNormalize_for_and_104_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_120_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_121_enex5 | NMP_ComputeSoftmaxNormalize_for_and_105_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_121_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_122_enex5 | NMP_ComputeSoftmaxNormalize_for_and_106_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_122_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_123_enex5 | NMP_ComputeSoftmaxNormalize_for_and_107_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_123_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_124_enex5 | NMP_ComputeSoftmaxNormalize_for_and_108_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_124_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_125_enex5 | NMP_ComputeSoftmaxNormalize_for_and_109_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_125_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_126_enex5 | NMP_ComputeSoftmaxNormalize_for_and_110_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_127_enex5 | NMP_ComputeSoftmaxNormalize_for_and_111_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_2_enexo <= NMP_ComputeSoftmaxNormalize_for_and_127_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_tmp
        | ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_2_enex5
        ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_acc_enexo
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_2_expret_qif_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_177_enex5 | NMP_ComputeRMSNormalize_for_and_161_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_177_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_178_enex5 | NMP_ComputeRMSNormalize_for_and_162_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_178_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_179_enex5 | NMP_ComputeRMSNormalize_for_and_163_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_179_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_180_enex5 | NMP_ComputeRMSNormalize_for_and_164_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_180_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_181_enex5 | NMP_ComputeRMSNormalize_for_and_165_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_181_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_182_enex5 | NMP_ComputeRMSNormalize_for_and_166_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_182_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_183_enex5 | NMP_ComputeRMSNormalize_for_and_167_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_183_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_184_enex5 | NMP_ComputeRMSNormalize_for_and_168_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_184_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_185_enex5 | NMP_ComputeRMSNormalize_for_and_169_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_185_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_186_enex5 | NMP_ComputeRMSNormalize_for_and_170_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_186_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_187_enex5 | NMP_ComputeRMSNormalize_for_and_171_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_187_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_188_enex5 | NMP_ComputeRMSNormalize_for_and_172_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_188_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_189_enex5 | NMP_ComputeRMSNormalize_for_and_173_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_189_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_190_enex5 | NMP_ComputeRMSNormalize_for_and_174_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_190_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_191_enex5 | NMP_ComputeRMSNormalize_for_and_175_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_191_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_192_enex5 | NMP_ComputeRMSNormalize_for_and_176_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_9_enexo <= NMP_ComputeRMSNormalize_for_and_192_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_cse |
        ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_4_enex5 ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_enexo
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_1_expret_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_15_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_106_enex5 | rva_out_reg_data_and_104_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_15_enexo <= rva_out_reg_data_and_106_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_15_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_107_enex5 | rva_out_reg_data_and_105_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_15_enexo <= rva_out_reg_data_and_107_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_sum_exp_39_4_sva_2_enexo <= 1'b1;
    end
    else if ( sum_exp_and_5_enex5 | sum_exp_and_4_enex5 ) begin
      reg_sum_exp_39_4_sva_2_enexo <= sum_exp_and_5_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_8_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_5_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_45_ssc | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_8_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_5_1_enexo <= NMP_PrepareWriteReq_and_45_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_5_1_enexo <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_9_enex5
        ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_5_1_enexo <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_1_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_87_enex5 | max_value_and_9_enex5 ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_1_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_87_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_1_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_86_enex5 | max_value_and_9_enex5 ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_1_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_86_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_1_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_88_enex5 | max_value_and_9_enex5 ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_1_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_88_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_max_value_26_0_sva_dfm_6_1_25_0_enexo <= 1'b1;
    end
    else if ( max_value_and_5_cse | max_value_and_9_enex5 ) begin
      reg_max_value_26_0_sva_dfm_6_1_25_0_enexo <= max_value_and_5_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_128_enex5 | NMP_ComputeSoftmaxNormalize_for_and_112_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_45_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_128_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_129_enex5 | NMP_ComputeSoftmaxNormalize_for_and_113_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_43_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_129_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_130_enex5 | NMP_ComputeSoftmaxNormalize_for_and_114_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_41_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_130_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_131_enex5 | NMP_ComputeSoftmaxNormalize_for_and_115_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_39_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_131_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_132_enex5 | NMP_ComputeSoftmaxNormalize_for_and_116_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_37_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_132_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_133_enex5 | NMP_ComputeSoftmaxNormalize_for_and_117_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_35_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_133_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_134_enex5 | NMP_ComputeSoftmaxNormalize_for_and_118_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_33_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_134_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_135_enex5 | NMP_ComputeSoftmaxNormalize_for_and_119_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_31_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_135_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_136_enex5 | NMP_ComputeSoftmaxNormalize_for_and_120_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_29_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_136_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_137_enex5 | NMP_ComputeSoftmaxNormalize_for_and_121_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_27_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_137_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_138_enex5 | NMP_ComputeSoftmaxNormalize_for_and_122_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_25_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_138_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_139_enex5 | NMP_ComputeSoftmaxNormalize_for_and_123_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_23_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_139_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_140_enex5 | NMP_ComputeSoftmaxNormalize_for_and_124_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_21_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_140_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_141_enex5 | NMP_ComputeSoftmaxNormalize_for_and_125_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_19_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_141_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_142_enex5 | NMP_ComputeSoftmaxNormalize_for_and_126_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_17_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_142_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxNormalize_for_and_143_enex5 | NMP_ComputeSoftmaxNormalize_for_and_127_enex5
        ) begin
      reg_NMP_ComputeSoftmaxNormalize_for_asn_itm_1_enexo <= NMP_ComputeSoftmaxNormalize_for_and_143_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_14_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_81_enex5 ) begin
      reg_input_fixed_14_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_13_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_82_enex5 ) begin
      reg_input_fixed_13_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_12_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_83_enex5 ) begin
      reg_input_fixed_12_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_11_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_84_enex5 ) begin
      reg_input_fixed_11_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_10_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_85_enex5 ) begin
      reg_input_fixed_10_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_9_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_86_enex5 ) begin
      reg_input_fixed_9_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_8_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_87_enex5 ) begin
      reg_input_fixed_8_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_7_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_88_enex5 ) begin
      reg_input_fixed_7_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_6_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_89_enex5 ) begin
      reg_input_fixed_6_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_5_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_90_enex5 ) begin
      reg_input_fixed_5_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_4_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_91_enex5 ) begin
      reg_input_fixed_4_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_3_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_ComputeSoftmaxExp_for_and_92_enex5 ) begin
      reg_input_fixed_3_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_96_enex5 | NMP_ComputeSoftmaxExp_for_and_93_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_96_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_97_enex5 | NMP_ComputeSoftmaxExp_for_and_94_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_16_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_97_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_98_enex5 | NMP_ComputeSoftmaxExp_for_and_95_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_itm_1_enexo <= NMP_ComputeSoftmaxExp_for_and_98_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_193_enex5 | NMP_ComputeRMSNormalize_for_and_177_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_193_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_194_enex5 | NMP_ComputeRMSNormalize_for_and_178_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_194_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_195_enex5 | NMP_ComputeRMSNormalize_for_and_179_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_195_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_196_enex5 | NMP_ComputeRMSNormalize_for_and_180_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_196_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_197_enex5 | NMP_ComputeRMSNormalize_for_and_181_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_197_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_198_enex5 | NMP_ComputeRMSNormalize_for_and_182_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_198_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_199_enex5 | NMP_ComputeRMSNormalize_for_and_183_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_199_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_200_enex5 | NMP_ComputeRMSNormalize_for_and_184_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_200_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_201_enex5 | NMP_ComputeRMSNormalize_for_and_185_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_201_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_202_enex5 | NMP_ComputeRMSNormalize_for_and_186_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_202_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_203_enex5 | NMP_ComputeRMSNormalize_for_and_187_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_203_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_204_enex5 | NMP_ComputeRMSNormalize_for_and_188_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_204_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_205_enex5 | NMP_ComputeRMSNormalize_for_and_189_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_205_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_206_enex5 | NMP_ComputeRMSNormalize_for_and_190_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_206_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_207_enex5 | NMP_ComputeRMSNormalize_for_and_191_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_207_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_208_enex5 | NMP_ComputeRMSNormalize_for_and_192_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_8_enexo <= NMP_ComputeRMSNormalize_for_and_208_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_13_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_63_enex5 | NMP_PrepareReadReq_and_56_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_1_itm_13_1_enexo <= NMP_PrepareReadReq_and_63_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_14_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_108_enex5 | rva_out_reg_data_and_106_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_14_enexo <= rva_out_reg_data_and_108_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_14_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_109_enex5 | rva_out_reg_data_and_107_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_14_enexo <= rva_out_reg_data_and_109_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_2_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_14_enex5
        | ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_13_enex5 ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_2_enexo
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_14_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_1_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_2_cse
        | operator_40_0_false_AC_TRN_AC_WRAP_1_and_enex5 ) begin
      reg_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_if_qr_lpi_1_dfm_st_1_1_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_qelse_and_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_sum_exp_39_4_sva_st_1_enexo_1 <= 1'b1;
    end
    else if ( sum_exp_and_3_enex5 | sum_exp_and_5_enex5 ) begin
      reg_sum_exp_39_4_sva_st_1_enexo_1 <= sum_exp_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_15_26_0_enexo <= 1'b1;
    end
    else if ( and_983_cse | NMP_RunFSM_switch_lp_and_342_enex5 ) begin
      reg_input_fixed_15_26_0_enexo <= and_983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_12_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_84_enex5 | NMP_PrepareWriteReq_and_63_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_12_enexo <= NMP_PrepareWriteReq_and_84_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_12_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_85_enex5 | NMP_PrepareWriteReq_and_64_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_12_1_enexo <= NMP_PrepareWriteReq_and_85_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_15_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_128_enex5 ) begin
      reg_exp_values_15_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_14_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_129_enex5 ) begin
      reg_exp_values_14_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_13_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_130_enex5 ) begin
      reg_exp_values_13_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_12_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_131_enex5 ) begin
      reg_exp_values_12_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_11_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_132_enex5 ) begin
      reg_exp_values_11_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_10_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_133_enex5 ) begin
      reg_exp_values_10_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_9_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_134_enex5 ) begin
      reg_exp_values_9_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_8_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_135_enex5 ) begin
      reg_exp_values_8_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_7_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_136_enex5 ) begin
      reg_exp_values_7_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_6_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_137_enex5 ) begin
      reg_exp_values_6_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_5_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_138_enex5 ) begin
      reg_exp_values_5_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_4_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_139_enex5 ) begin
      reg_exp_values_4_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_3_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_140_enex5 ) begin
      reg_exp_values_3_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_2_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_141_enex5 ) begin
      reg_exp_values_2_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_1_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_142_enex5 ) begin
      reg_exp_values_1_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_exp_values_0_enexo <= 1'b1;
    end
    else if ( and_1094_cse | NMP_ComputeSoftmaxNormalize_for_and_143_enex5 ) begin
      reg_exp_values_0_enexo <= and_1094_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_2_26_0_enexo <= 1'b1;
    end
    else if ( and_1067_cse | NMP_ComputeSoftmaxExp_for_and_96_enex5 ) begin
      reg_input_fixed_2_26_0_enexo <= and_1067_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_1_26_0_enexo <= 1'b1;
    end
    else if ( and_1067_cse | NMP_ComputeSoftmaxExp_for_and_97_enex5 ) begin
      reg_input_fixed_1_26_0_enexo <= and_1067_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_0_26_0_enexo <= 1'b1;
    end
    else if ( and_1067_cse | NMP_ComputeSoftmaxExp_for_and_98_enex5 ) begin
      reg_input_fixed_0_26_0_enexo <= and_1067_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_209_enex5 | NMP_ComputeRMSNormalize_for_and_193_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_209_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_210_enex5 | NMP_ComputeRMSNormalize_for_and_194_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_210_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_211_enex5 | NMP_ComputeRMSNormalize_for_and_195_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_211_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_212_enex5 | NMP_ComputeRMSNormalize_for_and_196_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_212_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_213_enex5 | NMP_ComputeRMSNormalize_for_and_197_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_213_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_214_enex5 | NMP_ComputeRMSNormalize_for_and_198_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_214_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_215_enex5 | NMP_ComputeRMSNormalize_for_and_199_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_215_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_216_enex5 | NMP_ComputeRMSNormalize_for_and_200_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_216_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_217_enex5 | NMP_ComputeRMSNormalize_for_and_201_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_217_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_218_enex5 | NMP_ComputeRMSNormalize_for_and_202_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_218_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_219_enex5 | NMP_ComputeRMSNormalize_for_and_203_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_219_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_220_enex5 | NMP_ComputeRMSNormalize_for_and_204_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_220_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_221_enex5 | NMP_ComputeRMSNormalize_for_and_205_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_221_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_222_enex5 | NMP_ComputeRMSNormalize_for_and_206_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_222_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_223_enex5 | NMP_ComputeRMSNormalize_for_and_207_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_223_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_224_enex5 | NMP_ComputeRMSNormalize_for_and_208_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_7_enexo <= NMP_ComputeRMSNormalize_for_and_224_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_12_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_76_enex5 | NMP_PrepareReadReq_and_57_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_12_1_enexo <= NMP_PrepareReadReq_and_76_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_13_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_110_enex5 | rva_out_reg_data_and_108_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_13_enexo <= rva_out_reg_data_and_110_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_13_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_111_enex5 | rva_out_reg_data_and_109_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_13_enexo <= rva_out_reg_data_and_111_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_9_cse |
        ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_14_enex5 ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1_enexo
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_9_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_fixed_1_26_0_enexo_1 <= 1'b1;
    end
    else if ( and_1067_cse | max_value_and_10_enex5 ) begin
      reg_input_fixed_1_26_0_enexo_1 <= and_1067_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_225_enex5 | NMP_ComputeRMSNormalize_for_and_209_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_225_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_226_enex5 | NMP_ComputeRMSNormalize_for_and_210_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_226_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_227_enex5 | NMP_ComputeRMSNormalize_for_and_211_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_227_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_228_enex5 | NMP_ComputeRMSNormalize_for_and_212_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_228_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_229_enex5 | NMP_ComputeRMSNormalize_for_and_213_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_229_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_230_enex5 | NMP_ComputeRMSNormalize_for_and_214_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_230_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_231_enex5 | NMP_ComputeRMSNormalize_for_and_215_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_231_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_232_enex5 | NMP_ComputeRMSNormalize_for_and_216_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_232_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_233_enex5 | NMP_ComputeRMSNormalize_for_and_217_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_233_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_234_enex5 | NMP_ComputeRMSNormalize_for_and_218_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_234_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_235_enex5 | NMP_ComputeRMSNormalize_for_and_219_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_235_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_236_enex5 | NMP_ComputeRMSNormalize_for_and_220_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_236_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_237_enex5 | NMP_ComputeRMSNormalize_for_and_221_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_237_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_238_enex5 | NMP_ComputeRMSNormalize_for_and_222_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_238_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_239_enex5 | NMP_ComputeRMSNormalize_for_and_223_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_239_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_240_enex5 | NMP_ComputeRMSNormalize_for_and_224_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_6_enexo <= NMP_ComputeRMSNormalize_for_and_240_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_12_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_112_enex5 | rva_out_reg_data_and_110_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_12_enexo <= rva_out_reg_data_and_112_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_12_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_113_enex5 | rva_out_reg_data_and_111_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_12_enexo <= rva_out_reg_data_and_113_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_241_enex5 | NMP_ComputeRMSNormalize_for_and_225_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_60_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_241_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_242_enex5 | NMP_ComputeRMSNormalize_for_and_226_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_242_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_243_enex5 | NMP_ComputeRMSNormalize_for_and_227_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_243_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_244_enex5 | NMP_ComputeRMSNormalize_for_and_228_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_244_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_245_enex5 | NMP_ComputeRMSNormalize_for_and_229_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_245_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_246_enex5 | NMP_ComputeRMSNormalize_for_and_230_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_246_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_247_enex5 | NMP_ComputeRMSNormalize_for_and_231_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_247_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_248_enex5 | NMP_ComputeRMSNormalize_for_and_232_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_248_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_249_enex5 | NMP_ComputeRMSNormalize_for_and_233_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_249_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_250_enex5 | NMP_ComputeRMSNormalize_for_and_234_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_250_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_251_enex5 | NMP_ComputeRMSNormalize_for_and_235_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_251_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_252_enex5 | NMP_ComputeRMSNormalize_for_and_236_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_252_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_253_enex5 | NMP_ComputeRMSNormalize_for_and_237_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_253_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_254_enex5 | NMP_ComputeRMSNormalize_for_and_238_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_254_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_255_enex5 | NMP_ComputeRMSNormalize_for_and_239_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_255_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_256_enex5 | NMP_ComputeRMSNormalize_for_and_240_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_5_enexo <= NMP_ComputeRMSNormalize_for_and_256_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_11_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_114_enex5 | rva_out_reg_data_and_112_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_11_enexo <= rva_out_reg_data_and_114_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_11_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_115_enex5 | rva_out_reg_data_and_113_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_11_enexo <= rva_out_reg_data_and_115_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_78_enex5 | NMP_PrepareWriteReq_and_65_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_9_enexo <= NMP_PrepareWriteReq_and_78_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_9_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_79_enex5 | NMP_PrepareWriteReq_and_66_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_9_1_enexo <= NMP_PrepareWriteReq_and_79_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_9_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_89_enex5 | NMP_PrepareWriteReq_and_67_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_9_2_enexo <= NMP_PrepareWriteReq_and_89_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_17 <= 1'b1;
    end
    else if ( NMP_RunFSM_switch_lp_and_126_enex5 | NMP_ComputeRMSNormalize_for_and_241_enex5
        ) begin
      reg_NMP_RunFSM_switch_lp_asn_104_itm_3_enexo_17 <= NMP_RunFSM_switch_lp_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_257_enex5 | NMP_ComputeRMSNormalize_for_and_242_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_58_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_257_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_258_enex5 | NMP_ComputeRMSNormalize_for_and_243_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_56_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_258_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_259_enex5 | NMP_ComputeRMSNormalize_for_and_244_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_54_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_259_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_260_enex5 | NMP_ComputeRMSNormalize_for_and_245_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_52_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_260_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_261_enex5 | NMP_ComputeRMSNormalize_for_and_246_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_50_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_261_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_262_enex5 | NMP_ComputeRMSNormalize_for_and_247_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_48_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_262_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_263_enex5 | NMP_ComputeRMSNormalize_for_and_248_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_46_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_263_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_264_enex5 | NMP_ComputeRMSNormalize_for_and_249_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_44_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_264_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_265_enex5 | NMP_ComputeRMSNormalize_for_and_250_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_42_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_265_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_266_enex5 | NMP_ComputeRMSNormalize_for_and_251_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_40_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_266_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_267_enex5 | NMP_ComputeRMSNormalize_for_and_252_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_38_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_267_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_268_enex5 | NMP_ComputeRMSNormalize_for_and_253_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_36_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_268_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_269_enex5 | NMP_ComputeRMSNormalize_for_and_254_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_269_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_270_enex5 | NMP_ComputeRMSNormalize_for_and_255_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_32_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_270_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_271_enex5 | NMP_ComputeRMSNormalize_for_and_256_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_4_enexo <= NMP_ComputeRMSNormalize_for_and_271_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_9_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_78_enex5 | NMP_PrepareReadReq_and_58_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_9_enexo <= NMP_PrepareReadReq_and_78_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_9_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_66_enex5 | NMP_PrepareReadReq_and_59_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_9_1_enexo <= NMP_PrepareReadReq_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_10_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_116_enex5 | rva_out_reg_data_and_114_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_10_enexo <= rva_out_reg_data_and_116_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_10_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_117_enex5 | rva_out_reg_data_and_115_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_10_enexo <= rva_out_reg_data_and_117_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo_2 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_67_enex5 | NMP_ComputeRMSNormalize_for_and_257_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_29_itm_2_enexo_2 <= NMP_ComputeSoftmaxExp_for_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo_2 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_68_enex5 | NMP_ComputeRMSNormalize_for_and_258_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_28_itm_2_enexo_2 <= NMP_ComputeSoftmaxExp_for_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo_2 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_69_enex5 | NMP_ComputeRMSNormalize_for_and_259_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_27_itm_2_enexo_2 <= NMP_ComputeSoftmaxExp_for_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo_2 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_70_enex5 | NMP_ComputeRMSNormalize_for_and_260_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_26_itm_2_enexo_2 <= NMP_ComputeSoftmaxExp_for_and_70_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo_2 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_21_enex5 | NMP_ComputeRMSNormalize_for_and_261_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_25_itm_2_enexo_2 <= NMP_ComputeSoftmaxExp_for_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_71_enex5 | NMP_ComputeRMSNormalize_for_and_262_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_24_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_71_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_72_enex5 | NMP_ComputeRMSNormalize_for_and_263_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_23_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_72_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_73_enex5 | NMP_ComputeRMSNormalize_for_and_264_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_22_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_73_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_74_enex5 | NMP_ComputeRMSNormalize_for_and_265_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_21_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_74_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_75_enex5 | NMP_ComputeRMSNormalize_for_and_266_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_20_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_75_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_76_enex5 | NMP_ComputeRMSNormalize_for_and_267_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_19_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_76_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_77_enex5 | NMP_ComputeRMSNormalize_for_and_268_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_18_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_77_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_272_enex5 | NMP_ComputeRMSNormalize_for_and_269_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_34_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_272_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSSqrtRecip_variance_and_1_ssc | NMP_ComputeRMSNormalize_for_and_270_enex5
        ) begin
      reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_1_enexo <= NMP_ComputeRMSSqrtRecip_variance_and_1_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSNormalize_for_and_273_enex5 | NMP_ComputeRMSNormalize_for_and_271_enex5
        ) begin
      reg_NMP_ComputeRMSNormalize_for_asn_itm_3_enexo <= NMP_ComputeRMSNormalize_for_and_273_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_9_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_118_enex5 | rva_out_reg_data_and_116_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_9_enexo <= rva_out_reg_data_and_118_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_9_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_119_enex5 | rva_out_reg_data_and_117_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_9_enexo <= rva_out_reg_data_and_119_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_93_enex5 | NMP_ComputeRMSNormalize_for_and_272_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_17_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_93_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeSoftmaxExp_for_and_95_enex5 | NMP_ComputeRMSNormalize_for_and_273_enex5
        ) begin
      reg_NMP_ComputeSoftmaxExp_for_asn_itm_2_enexo_1 <= NMP_ComputeSoftmaxExp_for_and_95_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_8_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_120_enex5 | rva_out_reg_data_and_118_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_8_enexo <= rva_out_reg_data_and_120_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_8_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_121_enex5 | rva_out_reg_data_and_119_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_8_enexo <= rva_out_reg_data_and_121_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_122_enex5 | rva_out_reg_data_and_120_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_7_enexo <= rva_out_reg_data_and_122_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_123_enex5 | rva_out_reg_data_and_121_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_7_enexo <= rva_out_reg_data_and_123_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_69_enex5 | NMP_PrepareWriteReq_and_68_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_5_enexo <= NMP_PrepareWriteReq_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_124_enex5 | rva_out_reg_data_and_122_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_6_enexo <= rva_out_reg_data_and_124_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_125_enex5 | rva_out_reg_data_and_123_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_6_enexo <= rva_out_reg_data_and_125_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_70_enex5 | NMP_PrepareWriteReq_and_69_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_4_enexo <= NMP_PrepareWriteReq_and_70_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_126_enex5 | rva_out_reg_data_and_124_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_5_enexo <= rva_out_reg_data_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_127_enex5 | rva_out_reg_data_and_125_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_5_enexo <= rva_out_reg_data_and_127_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_72_enex5 | NMP_PrepareWriteReq_and_70_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_3_enexo <= NMP_PrepareWriteReq_and_72_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_73_enex5 | NMP_PrepareWriteReq_and_71_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_3_enexo <= NMP_PrepareWriteReq_and_73_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_3_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_61_enex5 | NMP_PrepareReadReq_and_60_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_3_enexo <= NMP_PrepareReadReq_and_61_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_128_enex5 | rva_out_reg_data_and_126_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_4_enexo <= rva_out_reg_data_and_128_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_129_enex5 | rva_out_reg_data_and_127_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_4_enexo <= rva_out_reg_data_and_129_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_74_enex5 | NMP_PrepareWriteReq_and_72_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_2_enexo <= NMP_PrepareWriteReq_and_74_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_75_enex5 | NMP_PrepareWriteReq_and_73_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_2_enexo <= NMP_PrepareWriteReq_and_75_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_74_enex5 | NMP_PrepareReadReq_and_61_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_2_enexo_1 <= NMP_PrepareWriteReq_and_74_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_2_enexo_1 <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_75_enex5 | NMP_PrepareReadReq_and_62_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_2_enexo_1 <= NMP_PrepareWriteReq_and_75_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_130_enex5 | rva_out_reg_data_and_128_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_3_enexo <= rva_out_reg_data_and_130_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_131_enex5 | rva_out_reg_data_and_129_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_3_enexo <= rva_out_reg_data_and_131_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_76_enex5 | NMP_PrepareWriteReq_and_74_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_1_enexo <= NMP_PrepareWriteReq_and_76_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_77_enex5 | NMP_PrepareWriteReq_and_75_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_1_enexo <= NMP_PrepareWriteReq_and_77_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_132_enex5 | rva_out_reg_data_and_130_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_3_2_enexo <= rva_out_reg_data_and_132_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_133_enex5 | rva_out_reg_data_and_131_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_3_2_enexo <= rva_out_reg_data_and_133_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nmp_config_timestep_counter_enexo <= 1'b1;
    end
    else if ( and_1082_tmp | NMP_PrepareWriteReq_and_76_enex5 ) begin
      reg_nmp_config_timestep_counter_enexo <= and_1082_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nmp_config_vector_counter_enexo <= 1'b1;
    end
    else if ( and_1063_tmp | NMP_PrepareWriteReq_and_77_enex5 ) begin
      reg_nmp_config_vector_counter_enexo <= and_1063_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_132_enex5 ) begin
      reg_rva_out_reg_data_79_64_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_1_cse | rva_out_reg_data_and_133_enex5 ) begin
      reg_rva_out_reg_data_55_48_enexo <= rva_out_reg_data_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_1
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp |
        ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_enex5
        ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_1
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_1
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_3_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_1
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_1
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_3_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_1
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_1
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_3_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_1
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_2
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp |
        ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_3_enex5
        ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_2
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_2
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_4_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_2
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_2
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_4_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_2
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_2
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_4_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_2
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_3
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp |
        ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_4_enex5
        ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_3
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_3
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_5_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_1_enexo_3
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_4_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_3
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_5_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_24_12_sva_1_enexo_3
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_3
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_5_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_2_10_0_enexo_3
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_4
          <= 1'b1;
    end
    else if ( ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp |
        ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_m1_and_5_enex5
        ) begin
      reg_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_4_enexo_4
          <= ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mux_1_itm_2_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_9_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mux_1_itm_2_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_9_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1_enexo
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_8_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_10_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1_enexo
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_8_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1_enexo_1
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_8_enex5
        | ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_11_enex5
        ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_mul_psp_sva_1_enexo_1
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_8_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_12_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_64_enex5 | NMP_PrepareReadReq_and_63_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_1_itm_12_1_enexo <= NMP_PrepareReadReq_and_64_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_enexo <= 1'b1;
    end
    else if ( NMP_ComputeRMSSqrtRecip_variance_and_1_ssc | NMP_ComputeRMSSqrtRecip_variance_and_enex5
        ) begin
      reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_enexo <= NMP_ComputeRMSSqrtRecip_variance_and_1_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_1_enexo_1 <= 1'b1;
    end
    else if ( NMP_ComputeRMSSqrtRecip_variance_and_1_ssc | NMP_ComputeRMSSqrtRecip_variance_and_2_enex5
        ) begin
      reg_NMP_ComputeRMSSqrtRecip_variance_acc_psp_sva_1_1_enexo_1 <= NMP_ComputeRMSSqrtRecip_variance_and_1_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_11_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_65_enex5 | NMP_PrepareReadReq_and_64_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_1_itm_11_1_enexo <= NMP_PrepareReadReq_and_65_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_10_1_enexo <= 1'b1;
    end
    else if ( NMPRun_wen | NMP_PrepareReadReq_and_65_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_10_1_enexo <= NMPRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_80_enex5 | NMP_PrepareWriteReq_and_78_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_8_enexo <= NMP_PrepareWriteReq_and_80_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_8_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_81_enex5 | NMP_PrepareWriteReq_and_79_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_8_1_enexo <= NMP_PrepareWriteReq_and_81_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_8_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_67_enex5 | NMP_PrepareReadReq_and_66_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_8_1_enexo <= NMP_PrepareReadReq_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_82_enex5 | NMP_PrepareWriteReq_and_80_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_7_enexo <= NMP_PrepareWriteReq_and_82_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_7_1_enexo <= 1'b1;
    end
    else if ( ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_36_ssc
        | NMP_PrepareWriteReq_and_81_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_7_1_enexo <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_36_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_7_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_40_ssc | NMP_PrepareReadReq_and_67_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_7_1_enexo <= NMP_PrepareReadReq_and_40_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_68_enex5 | NMP_PrepareWriteReq_and_82_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_6_enexo <= NMP_PrepareWriteReq_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_6_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_69_enex5 | NMP_PrepareReadReq_and_68_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_6_enexo <= NMP_PrepareReadReq_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_5_1_enexo_1 <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_45_ssc | NMP_PrepareWriteReq_and_83_enex5 )
        begin
      reg_NMP_PrepareWriteReq_asn_1_itm_5_1_enexo_1 <= NMP_PrepareWriteReq_and_45_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_5_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_72_enex5 | NMP_PrepareReadReq_and_69_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_5_enexo <= NMP_PrepareReadReq_and_72_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_5_1_enexo_1 <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc
        | NMP_PrepareReadReq_and_70_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_5_1_enexo_1 <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_2_enexo_1
          <= 1'b1;
    end
    else if ( ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc
        | NMP_PrepareReadReq_and_71_enex5 ) begin
      reg_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_slc_ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_38_25_11_0_itm_1_2_enexo_1
          <= ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_input_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_4_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_60_enex5 | NMP_PrepareReadReq_and_72_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_4_enexo <= NMP_PrepareReadReq_and_60_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_15_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_74_enex5 | NMP_PrepareReadReq_and_73_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_1_itm_15_1_enexo <= NMP_PrepareReadReq_and_74_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_14_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_56_enex5 | NMP_PrepareReadReq_and_74_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_1_itm_14_1_enexo <= NMP_PrepareReadReq_and_56_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_11_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_87_enex5 | NMP_PrepareWriteReq_and_84_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_11_enexo <= NMP_PrepareWriteReq_and_87_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_11_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_88_enex5 | NMP_PrepareWriteReq_and_85_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_11_1_enexo <= NMP_PrepareWriteReq_and_88_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_11_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_96_enex5 | NMP_PrepareWriteReq_and_86_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_11_2_enexo <= NMP_PrepareWriteReq_and_96_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_11_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_85_enex5 | NMP_PrepareReadReq_and_75_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_11_enexo <= NMP_PrepareReadReq_and_85_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_11_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_77_enex5 | NMP_PrepareReadReq_and_76_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_11_1_enexo <= NMP_PrepareReadReq_and_77_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_10_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_65_enex5 | NMP_PrepareWriteReq_and_87_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_10_enexo <= NMP_PrepareWriteReq_and_65_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_10_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_66_enex5 | NMP_PrepareWriteReq_and_88_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_10_1_enexo <= NMP_PrepareWriteReq_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_59_enex5 | NMP_PrepareReadReq_and_77_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_1_enexo <= NMP_PrepareReadReq_and_59_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_8_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_90_enex5 | NMP_PrepareWriteReq_and_89_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_8_2_enexo <= NMP_PrepareWriteReq_and_90_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_8_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_80_enex5 | NMP_PrepareReadReq_and_78_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_8_enexo <= NMP_PrepareReadReq_and_80_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_8_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_81_enex5 | NMP_PrepareReadReq_and_79_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_1_itm_8_2_enexo <= NMP_PrepareReadReq_and_81_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_7_2_enexo <= 1'b1;
    end
    else if ( ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_36_ssc
        | NMP_PrepareWriteReq_and_90_enex5 ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_7_2_enexo <= ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_36_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_7_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_68_enex5 | NMP_PrepareReadReq_and_80_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_7_enexo <= NMP_PrepareReadReq_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_7_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_40_ssc | NMP_PrepareReadReq_and_81_enex5 ) begin
      reg_NMP_PrepareReadReq_asn_1_itm_7_2_enexo <= NMP_PrepareReadReq_and_40_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_14_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_94_enex5 | NMP_PrepareWriteReq_and_91_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_14_enexo <= NMP_PrepareWriteReq_and_94_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_14_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_95_enex5 | NMP_PrepareWriteReq_and_92_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_14_1_enexo <= NMP_PrepareWriteReq_and_95_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_14_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_98_enex5 | NMP_PrepareWriteReq_and_93_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_14_2_enexo <= NMP_PrepareWriteReq_and_98_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_14_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_87_enex5 | NMP_PrepareReadReq_and_82_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_14_enexo <= NMP_PrepareReadReq_and_87_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_14_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_84_enex5 | NMP_PrepareReadReq_and_83_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_14_1_enexo <= NMP_PrepareReadReq_and_84_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_13_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_63_enex5 | NMP_PrepareWriteReq_and_94_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_13_enexo <= NMP_PrepareWriteReq_and_63_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_13_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_64_enex5 | NMP_PrepareWriteReq_and_95_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_2_itm_13_1_enexo <= NMP_PrepareWriteReq_and_64_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_13_1_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_57_enex5 | NMP_PrepareReadReq_and_84_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_13_1_enexo <= NMP_PrepareReadReq_and_57_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_10_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_67_enex5 | NMP_PrepareWriteReq_and_96_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_10_2_enexo <= NMP_PrepareWriteReq_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_58_enex5 | NMP_PrepareReadReq_and_85_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_10_enexo <= NMP_PrepareReadReq_and_58_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_12_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_86_enex5 | NMP_PrepareWriteReq_and_97_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_12_2_enexo <= NMP_PrepareWriteReq_and_86_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_12_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_75_enex5 | NMP_PrepareReadReq_and_86_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_12_enexo <= NMP_PrepareReadReq_and_75_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_13_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_97_enex5 | NMP_PrepareWriteReq_and_98_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_13_2_enexo <= NMP_PrepareWriteReq_and_97_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_13_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_86_enex5 | NMP_PrepareReadReq_and_87_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_13_enexo <= NMP_PrepareReadReq_and_86_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareReadReq_asn_2_itm_15_enexo <= 1'b1;
    end
    else if ( NMP_PrepareReadReq_and_82_enex5 | NMP_PrepareReadReq_and_88_enex5 )
        begin
      reg_NMP_PrepareReadReq_asn_2_itm_15_enexo <= NMP_PrepareReadReq_and_82_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_15_2_enexo <= 1'b1;
    end
    else if ( NMP_PrepareWriteReq_and_93_enex5 | NMP_PrepareWriteReq_and_99_enex5
        ) begin
      reg_NMP_PrepareWriteReq_asn_1_itm_15_2_enexo <= NMP_PrepareWriteReq_and_93_enex5;
    end
  end
  assign NMP_PrepareReadReq_or_nl = ((~ NMP_RunFSM_switch_lp_conc_itm_10_2) & xor_3_ssc)
      | (NMP_RunFSM_switch_lp_conc_itm_10_2 & xor_3_ssc);
  assign nl_NMP_ConvertOutputToAdpfloat_for_16_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_1_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_16_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_16_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_15_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_1_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_16_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_1_sva_1_6);
  assign operator_5_true_not_127_nl = ~ NMP_ConvertOutputToAdpfloat_for_16_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_16_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_15_nl,
      4'b1111, operator_5_true_not_127_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_1_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_16_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_15_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_1_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_16_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_1_sva_1_6);
  assign operator_5_true_1_not_127_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_16_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_16_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_15_nl,
      4'b1111, operator_5_true_1_not_127_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_15_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_17_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_15_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_15_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_14_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_17_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_15_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_17_sva_1_6);
  assign operator_5_true_not_126_nl = ~ NMP_ConvertOutputToAdpfloat_for_15_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_17_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_14_nl,
      4'b1111, operator_5_true_not_126_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_17_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_15_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_14_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_17_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_15_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_17_sva_1_6);
  assign operator_5_true_1_not_126_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_15_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_17_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_14_nl,
      4'b1111, operator_5_true_1_not_126_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_14_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_16_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_14_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_14_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_13_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_16_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_14_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_16_sva_1_6);
  assign operator_5_true_not_125_nl = ~ NMP_ConvertOutputToAdpfloat_for_14_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_18_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_13_nl,
      4'b1111, operator_5_true_not_125_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_16_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_14_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_13_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_16_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_14_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_16_sva_1_6);
  assign operator_5_true_1_not_125_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_14_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_18_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_13_nl,
      4'b1111, operator_5_true_1_not_125_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_13_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_15_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_13_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_13_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_12_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_15_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_13_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_15_sva_1_6);
  assign operator_5_true_not_124_nl = ~ NMP_ConvertOutputToAdpfloat_for_13_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_19_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_12_nl,
      4'b1111, operator_5_true_not_124_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_15_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_13_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_12_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_15_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_13_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_15_sva_1_6);
  assign operator_5_true_1_not_124_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_13_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_19_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_12_nl,
      4'b1111, operator_5_true_1_not_124_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_12_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_14_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_12_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_12_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_11_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_14_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_12_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_14_sva_1_6);
  assign operator_5_true_not_123_nl = ~ NMP_ConvertOutputToAdpfloat_for_12_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_20_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_11_nl,
      4'b1111, operator_5_true_not_123_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_14_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_12_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_11_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_14_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_12_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_14_sva_1_6);
  assign operator_5_true_1_not_123_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_12_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_20_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_11_nl,
      4'b1111, operator_5_true_1_not_123_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_11_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_13_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_11_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_11_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_10_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_13_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_11_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_13_sva_1_6);
  assign operator_5_true_not_122_nl = ~ NMP_ConvertOutputToAdpfloat_for_11_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_21_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_10_nl,
      4'b1111, operator_5_true_not_122_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_13_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_11_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_10_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_13_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_11_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_13_sva_1_6);
  assign operator_5_true_1_not_122_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_11_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_21_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_10_nl,
      4'b1111, operator_5_true_1_not_122_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_10_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_12_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_10_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_10_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_9_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_12_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_10_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_12_sva_1_6);
  assign operator_5_true_not_121_nl = ~ NMP_ConvertOutputToAdpfloat_for_10_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_22_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_9_nl,
      4'b1111, operator_5_true_not_121_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_12_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_10_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_9_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_12_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_10_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_12_sva_1_6);
  assign operator_5_true_1_not_121_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_10_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_22_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_9_nl,
      4'b1111, operator_5_true_1_not_121_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_9_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_11_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_9_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_9_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_8_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_11_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_9_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_11_sva_1_6);
  assign operator_5_true_not_120_nl = ~ NMP_ConvertOutputToAdpfloat_for_9_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_23_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_8_nl,
      4'b1111, operator_5_true_not_120_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_11_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_9_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_8_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_11_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_9_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_11_sva_1_6);
  assign operator_5_true_1_not_120_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_9_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_23_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_8_nl,
      4'b1111, operator_5_true_1_not_120_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_8_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_10_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_8_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_8_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_7_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_10_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_8_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_10_sva_1_6);
  assign operator_5_true_not_119_nl = ~ NMP_ConvertOutputToAdpfloat_for_8_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_24_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_7_nl,
      4'b1111, operator_5_true_not_119_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_10_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_8_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_7_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_10_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_8_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_10_sva_1_6);
  assign operator_5_true_1_not_119_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_8_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_24_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_7_nl,
      4'b1111, operator_5_true_1_not_119_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_7_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_9_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_7_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_7_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_6_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_9_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_7_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_9_sva_1_6);
  assign operator_5_true_not_118_nl = ~ NMP_ConvertOutputToAdpfloat_for_7_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_25_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_6_nl,
      4'b1111, operator_5_true_not_118_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_9_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_7_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_6_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_9_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_7_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_9_sva_1_6);
  assign operator_5_true_1_not_118_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_7_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_25_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_6_nl,
      4'b1111, operator_5_true_1_not_118_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_6_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_8_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_6_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_6_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_5_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_8_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_6_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_8_sva_1_6);
  assign operator_5_true_not_117_nl = ~ NMP_ConvertOutputToAdpfloat_for_6_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_26_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_5_nl,
      4'b1111, operator_5_true_not_117_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_8_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_6_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_5_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_8_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_6_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_8_sva_1_6);
  assign operator_5_true_1_not_117_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_6_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_26_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_5_nl,
      4'b1111, operator_5_true_1_not_117_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_5_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_7_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_5_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_5_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_4_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_7_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_5_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_7_sva_1_6);
  assign operator_5_true_not_116_nl = ~ NMP_ConvertOutputToAdpfloat_for_5_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_27_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_4_nl,
      4'b1111, operator_5_true_not_116_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_7_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_5_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_4_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_7_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_5_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_7_sva_1_6);
  assign operator_5_true_1_not_116_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_5_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_27_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_4_nl,
      4'b1111, operator_5_true_1_not_116_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_4_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_6_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_4_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_4_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_3_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_6_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_4_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_6_sva_1_6);
  assign operator_5_true_not_115_nl = ~ NMP_ConvertOutputToAdpfloat_for_4_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_28_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_3_nl,
      4'b1111, operator_5_true_not_115_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_6_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_4_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_3_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_6_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_4_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_6_sva_1_6);
  assign operator_5_true_1_not_115_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_4_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_28_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_3_nl,
      4'b1111, operator_5_true_1_not_115_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_3_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_5_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_3_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_3_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_2_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_5_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_3_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_5_sva_1_6);
  assign operator_5_true_not_114_nl = ~ NMP_ConvertOutputToAdpfloat_for_3_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_29_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_2_nl,
      4'b1111, operator_5_true_not_114_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_5_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_3_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_2_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_5_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_3_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_5_sva_1_6);
  assign operator_5_true_1_not_114_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_3_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_29_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_2_nl,
      4'b1111, operator_5_true_1_not_114_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_2_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_4_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_2_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_2_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_1_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_4_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_2_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_4_sva_1_6);
  assign operator_5_true_not_113_nl = ~ NMP_ConvertOutputToAdpfloat_for_2_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_30_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_1_nl,
      4'b1111, operator_5_true_not_113_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_4_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_2_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_1_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_4_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_2_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_4_sva_1_6);
  assign operator_5_true_1_not_113_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_2_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_30_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_1_nl,
      4'b1111, operator_5_true_1_not_113_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_1_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      =  -out_float_round_32_if_m_1_3_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_for_1_out_adp_set_value_ac_float_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_1_out_adp_set_value_ac_float_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_else_1_else_mux_nl = MUX_v_4_2_2(out_float_round_32_if_m_1_3_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_for_1_out_adp_set_value_ac_float_else_1_else_if_acc_nl,
      out_float_round_32_if_m_1_3_sva_1_6);
  assign operator_5_true_not_112_nl = ~ NMP_ConvertOutputToAdpfloat_for_1_operator_5_true_slc_operator_5_true_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_nor_31_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_else_1_else_mux_nl,
      4'b1111, operator_5_true_not_112_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      =  -out_float_round_32_1_if_m_1_3_sva_1_3_0;
  assign NMP_ConvertOutputToAdpfloat_1_for_1_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl[3:0];
  assign out_adp_set_value_ac_float_1_else_1_else_mux_nl = MUX_v_4_2_2(out_float_round_32_1_if_m_1_3_sva_1_3_0,
      NMP_ConvertOutputToAdpfloat_1_for_1_out_adp_set_value_ac_float_1_else_1_else_if_acc_nl,
      out_float_round_32_1_if_m_1_3_sva_1_6);
  assign operator_5_true_1_not_112_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_1_operator_5_true_1_slc_operator_5_true_1_acc_2_svs_mx0w0;
  assign out_adp_set_value_ac_float_1_nor_31_nl = ~(MUX_v_4_2_2(out_adp_set_value_ac_float_1_else_1_else_mux_nl,
      4'b1111, operator_5_true_1_not_112_nl));
  assign nl_NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_30_nl = ~ NMP_ConvertOutputToAdpfloat_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_15_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_29_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_29_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_15_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_29_nl = ~ NMP_ConvertOutputToAdpfloat_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_14_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_27_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_27_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_14_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_28_nl = ~ NMP_ConvertOutputToAdpfloat_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_13_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_13_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_27_nl = ~ NMP_ConvertOutputToAdpfloat_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_12_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_23_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_23_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_12_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_26_nl = ~ NMP_ConvertOutputToAdpfloat_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_11_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_21_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_21_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_11_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_25_nl = ~ NMP_ConvertOutputToAdpfloat_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_10_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_19_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_19_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_10_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_24_nl = ~ NMP_ConvertOutputToAdpfloat_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_9_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_17_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_17_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_9_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_23_nl = ~ NMP_ConvertOutputToAdpfloat_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_8_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_15_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_15_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_8_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_22_nl = ~ NMP_ConvertOutputToAdpfloat_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_7_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_7_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_21_nl = ~ NMP_ConvertOutputToAdpfloat_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_6_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_11_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_11_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_6_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_20_nl = ~ NMP_ConvertOutputToAdpfloat_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_5_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_9_nl =
      MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_9_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_5_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_19_nl = ~ NMP_ConvertOutputToAdpfloat_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_4_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_7_nl =
      MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_7_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_4_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_18_nl = ~ NMP_ConvertOutputToAdpfloat_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_3_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_5_nl =
      MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_5_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_3_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_17_nl = ~ NMP_ConvertOutputToAdpfloat_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_2_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_3_nl =
      MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_3_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_2_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_16_nl = ~ NMP_ConvertOutputToAdpfloat_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_ls_4_0_1_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl =
      MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl +
      conv_u2s_1_5(out_float_round_32_rnd_ovfl_1_sva_1);
  assign NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_not_nl = ~ NMP_ConvertOutputToAdpfloat_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_31_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_31_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_30_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_16_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_15_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_29_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_29_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_15_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_29_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_15_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_14_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_27_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_27_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_14_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_28_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_14_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_13_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_25_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_25_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_13_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_27_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_13_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_12_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_23_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_23_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_12_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_26_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_12_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_11_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_21_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_21_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_11_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_25_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_11_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_10_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_19_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_19_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_10_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_24_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_10_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_9_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_17_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_17_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_9_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_23_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_9_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_8_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_15_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_15_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_8_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_22_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_8_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_7_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_13_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_13_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_7_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_21_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_7_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_6_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_11_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_11_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_6_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_20_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_6_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_5_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_9_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_9_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_5_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_19_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_5_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_4_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_7_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_7_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_4_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_18_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_4_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_3_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_5_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_5_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_3_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_17_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_3_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_2_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_3_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_3_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_2_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_16_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_2_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = (~ out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_ls_4_0_1_sva_1) + 5'b01011;
  assign NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_1_nl
      = MUX_v_5_2_2(5'b10000, NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_slc_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_4_svs_st_1);
  assign nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_1_nl
      + conv_u2s_1_5(out_float_round_32_1_rnd_ovfl_1_sva_1);
  assign NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl
      = nl_NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_qelse_acc_nl[4:0];
  assign out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_not_nl = ~ NMP_ConvertOutputToAdpfloat_1_for_1_out_float_assign_from_0_0_32_12_AC_TRN_AC_WRAP_1_if_and_svs_st_1;
  assign nl_NMP_ComputeSoftmaxExp_for_16_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_30_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_15_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_29_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_14_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_28_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_13_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_27_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_12_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_26_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_11_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_25_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_10_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_24_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_9_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_23_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_8_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_22_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_7_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_21_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_6_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_20_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_5_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_19_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_4_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_18_itm_2)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_3_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_17_itm_3)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_2_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_16_itm_3)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign nl_NMP_ComputeSoftmaxExp_for_1_acc_1_itm_1  = conv_s2s_27_28(NMP_ComputeSoftmaxExp_for_asn_itm_3)
      + conv_s2s_27_28({(~ max_value_mux_1_itm) , (~ max_value_mux_2_itm)}) + 28'b0000000000000000000000000001;
  assign NMP_RunFSM_switch_lp_not_64_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_51_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_16_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_64_nl);
  assign NMP_RunFSM_switch_lp_not_65_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_50_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_15_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_65_nl);
  assign NMP_RunFSM_switch_lp_not_66_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_49_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_14_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_66_nl);
  assign NMP_RunFSM_switch_lp_not_67_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_48_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_13_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_67_nl);
  assign NMP_RunFSM_switch_lp_not_68_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_47_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_12_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_68_nl);
  assign NMP_RunFSM_switch_lp_not_69_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_46_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_11_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_69_nl);
  assign NMP_RunFSM_switch_lp_not_70_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_45_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_10_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_70_nl);
  assign NMP_RunFSM_switch_lp_not_71_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_44_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_9_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_71_nl);
  assign NMP_RunFSM_switch_lp_not_72_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_43_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_8_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_72_nl);
  assign NMP_RunFSM_switch_lp_not_73_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_42_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_7_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_73_nl);
  assign NMP_RunFSM_switch_lp_not_74_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_41_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_6_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_74_nl);
  assign NMP_RunFSM_switch_lp_not_75_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_40_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_5_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_75_nl);
  assign NMP_RunFSM_switch_lp_not_76_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_NMP_RunFSM_switch_lp_and_39_nl = MUX_v_27_2_2(27'b000000000000000000000000000,
      NMP_ConvertInputToFixed_for_4_in_float_to_ac_fixed_lshift_1_itm, NMP_RunFSM_switch_lp_not_76_nl);
  assign mux_277_nl = MUX_s_1_2_2(is_start_sva, and_1236_itm, start_PopNB_mioi_return_rsc_z_mxwt);
  assign NMP_RunFSM_switch_lp_or_41_nl = NMP_RunFSM_switch_lp_equal_tmp_22 | NMP_RunFSM_switch_lp_equal_tmp_18_1
      | NMP_RunFSM_switch_lp_equal_tmp_20 | NMP_RunFSM_switch_lp_equal_tmp_23 | NMP_RunFSM_switch_lp_equal_tmp_17
      | NMP_RunFSM_switch_lp_equal_tmp_19 | NMP_RunFSM_switch_lp_equal_tmp_21 | NMP_RunFSM_switch_lp_equal_tmp_24
      | NMP_RunFSM_switch_lp_equal_tmp_25 | NMP_RunFSM_switch_lp_equal_tmp_11_1 |
      NMP_RunFSM_switch_lp_equal_tmp_12_1 | NMP_RunFSM_switch_lp_or_tmp_1;
  assign NMP_RunFSM_switch_lp_mux_32_nl = MUX_s_1_2_2(mux_277_nl, is_start_sva, NMP_RunFSM_switch_lp_or_41_nl);
  assign NMP_RunFSM_switch_lp_not_77_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_not_78_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign NMP_RunFSM_switch_lp_not_51_nl = ~ NMP_RunFSM_switch_lp_equal_tmp_1;
  assign nl_operator_16_false_acc_2_nl = nmp_config_timestep_counter_sva + 16'b0000000000000001;
  assign operator_16_false_acc_2_nl = nl_operator_16_false_acc_2_nl[15:0];
  assign mux_222_nl = MUX_s_1_2_2((~ mux_cse), operator_16_false_acc_2_itm_17, NMP_RunFSM_switch_lp_and_2_rgt);
  assign nl_nmp_config_vector_counter_sva_3_1  = nmp_config_vector_counter_sva_mx1
      + 8'b00000001;
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_psp_sva
      = conv_s2u_9_11(ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_mx0w0[18:10])
      + ({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_40_16_true_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_itm});
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_acc_itm
      = conv_s2u_9_11(ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10])
      + ({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_40_16_false_AC_TRN_AC_WRAP_40_16_true_AC_TRN_AC_WRAP_output_pwl_mux_1_itm});
  assign mux_171_nl = MUX_s_1_2_2(mux_tmp_151, mux_tmp_161, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_167_nl = MUX_s_1_2_2(mux_tmp_147, mux_146_cse, large_rsp_PopNB_mioi_return_rsc_z_mxwt);
  assign mux_168_nl = MUX_s_1_2_2(mux_149_itm, mux_167_nl, NMP_RunFSM_switch_lp_equal_tmp_11_1);
  assign mux_166_nl = MUX_s_1_2_2(mux_219_cse, mux_146_cse, NMP_RunFSM_switch_lp_and_8_cse_1);
  assign mux_169_nl = MUX_s_1_2_2(mux_168_nl, mux_166_nl, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign or_836_nl = (~((~ NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2) |
      NMP_RunFSM_switch_lp_or_73_tmp)) | NMP_UpdateFSM_switch_lp_equal_tmp_1 | NMP_UpdateFSM_switch_lp_nor_tmp_1;
  assign mux_162_nl = MUX_s_1_2_2(mux_tmp_142, nor_tmp_19, or_836_nl);
  assign mux_163_nl = MUX_s_1_2_2(mux_tmp_156, mux_162_nl, NMP_RunFSM_switch_lp_and_8_cse_1);
  assign mux_164_nl = MUX_s_1_2_2(mux_163_nl, mux_tmp_161, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign mux_170_nl = MUX_s_1_2_2(mux_169_nl, mux_164_nl, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_172_nl = MUX_s_1_2_2(mux_171_nl, mux_170_nl, state_1_sva);
  assign mux_173_nl = MUX_s_1_2_2(mux_172_nl, mux_tmp_152, state_0_sva);
  assign mux_157_nl = MUX_s_1_2_2(mux_tmp_150, nor_tmp_19, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign mux_158_nl = MUX_s_1_2_2(mux_157_nl, mux_tmp_156, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_282_nl = MUX_s_1_2_2(mux_tmp_142, nor_tmp_19, or_tmp_129);
  assign and_894_nl = NMP_RunFSM_switch_lp_equal_tmp_11_1 & NMP_UpdateFSM_case_0_if_1_ac_int_cctor_lpi_1_dfm_2;
  assign mux_153_nl = MUX_s_1_2_2(mux_282_nl, nor_tmp_19, and_894_nl);
  assign mux_154_nl = MUX_s_1_2_2(mux_tmp_150, mux_153_nl, NMP_RunFSM_switch_lp_equal_tmp_12_1);
  assign mux_155_nl = MUX_s_1_2_2(mux_154_nl, mux_tmp_143, NMP_RunFSM_switch_lp_equal_tmp_1);
  assign mux_159_nl = MUX_s_1_2_2(mux_158_nl, mux_155_nl, or_801_cse);
  assign mux_160_nl = MUX_s_1_2_2(mux_tmp_152, mux_159_nl, nor_tmp_17);
  assign mux_174_nl = MUX_s_1_2_2(mux_173_nl, mux_160_nl, state_3_sva);
  assign mux_175_nl = MUX_s_1_2_2((~ mux_174_nl), mux_tmp_139, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_176_nl = MUX_s_1_2_2(mux_tmp_140, mux_175_nl, while_stage_0_3);
  assign or_830_nl = (~ while_stage_0_3) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ mux_tmp_152);
  assign mux_177_nl = MUX_s_1_2_2(mux_176_nl, or_830_nl, state_2_sva);
  assign nand_2_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & (~ mux_tmp_139));
  assign mux_141_nl = MUX_s_1_2_2(mux_tmp_140, nand_2_nl, while_stage_0_3);
  assign or_820_nl = state_2_sva | mux_141_nl;
  assign or_815_nl = NMP_UpdateFSM_switch_lp_equal_tmp_2_1 | NMP_UpdateFSM_switch_lp_equal_tmp_3_1
      | NMP_UpdateFSM_switch_lp_equal_tmp_5_1 | NMP_UpdateFSM_switch_lp_equal_tmp_6_1;
  assign mux_178_nl = MUX_s_1_2_2(mux_177_nl, or_820_nl, or_815_nl);
  assign and_671_nl = (~ mux_178_nl) & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign nl_NMP_ComputeSoftmaxSum_for_acc_7_itm_1  = conv_u2u_32_34(exp_values_5_sva_mx1)
      + conv_u2u_32_34(exp_values_4_sva_mx1) + conv_u2u_32_34(exp_values_3_sva_mx1);
  assign nl_NMP_ComputeSoftmaxSum_for_acc_8_itm_1  = conv_u2u_32_34(exp_values_7_sva_mx1)
      + conv_u2u_32_34(exp_values_8_sva_mx1) + conv_u2u_32_34(exp_values_6_sva_mx1);
  assign nl_NMP_ComputeSoftmaxSum_for_acc_9_itm_1  = conv_u2u_32_34(exp_values_9_sva_mx1)
      + conv_u2u_32_34(exp_values_10_sva_mx1) + conv_u2u_32_34(exp_values_11_sva_mx1);
  assign nl_NMP_ComputeSoftmaxSum_for_acc_11_itm_1  = conv_u2u_32_34(exp_values_2_sva_mx1)
      + conv_u2u_32_34(exp_values_1_sva_mx1) + conv_u2u_32_34(exp_values_0_sva_mx1);
  assign nl_NMP_ComputeSoftmaxSum_for_acc_12_itm_1  = conv_u2u_32_33(exp_values_12_sva_mx1)
      + conv_u2u_32_33(exp_values_13_sva_mx1);
  assign nl_NMP_ComputeSoftmaxSum_for_acc_13_itm_1  = conv_u2u_32_33(exp_values_14_sva_mx1)
      + conv_u2u_32_33(exp_values_15_sva_mx1);
  assign nl_ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_qr_6_0_sva_1 
      = ({1'b1 , (~ leading_sign_40_0_out_1)}) + 7'b0010001;
  assign nl_NMP_ComputeRMSSumSq_for_acc_3_nl = conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_z[53:16]);
  assign NMP_ComputeRMSSumSq_for_acc_3_nl = nl_NMP_ComputeRMSSumSq_for_acc_3_nl[39:0];
  assign nl_NMP_ComputeRMSSumSq_for_acc_nl = NMP_ComputeRMSSumSq_for_acc_3_nl + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_z[53:16])
      + conv_s2s_38_40(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_z[53:16]);
  assign NMP_ComputeRMSSumSq_for_acc_nl = nl_NMP_ComputeRMSSumSq_for_acc_nl[39:0];
  assign nmp_config_ConfigRead_not_12_nl = ~ nmp_config_ConfigRead_unequal_tmp_1;
  assign nmp_config_ConfigRead_not_10_nl = ~ nmp_config_ConfigRead_unequal_tmp_1;
  assign nmp_config_ConfigRead_not_9_nl = ~ nmp_config_ConfigRead_unequal_tmp_1;
  assign nmp_config_ConfigRead_not_6_nl = ~ nmp_config_ConfigRead_unequal_tmp_1;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_nl
      = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[33:32]==2'b00)
      & NMP_RunFSM_switch_lp_conc_itm_7_1;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_1_nl
      = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[33:32]==2'b01)
      & NMP_RunFSM_switch_lp_conc_itm_7_1;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_2_nl
      = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[33:32]==2'b10)
      & NMP_RunFSM_switch_lp_conc_itm_7_1;
  assign ac_math_ac_sqrt_pwl_AC_TRN_40_16_AC_TRN_AC_WRAP_40_16_AC_TRN_AC_WRAP_normalized_output_and_3_nl
      = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z[33:32]==2'b11)
      & NMP_RunFSM_switch_lp_conc_itm_7_1;
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux_nl
      = MUX_s_1_2_2(out_adp_set_value_ac_float_1_asn_15_itm_6_rsp_0, out_adp_set_value_ac_float_asn_15_itm_6_rsp_0,
      and_835_itm);
  assign and_833_nl = NMP_RunFSM_switch_lp_conc_itm_7_3 & (~ NMP_RunFSM_switch_lp_conc_itm_7_1);
  assign and_836_nl = and_dcpl_832 & (~ NMP_RunFSM_switch_lp_conc_itm_7_2);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux1h_60_nl
      = MUX1HOT_v_2_5_2(2'b01, 2'b10, out_adp_set_value_ac_float_1_asn_15_itm_6_rsp_1,
      out_adp_set_value_ac_float_asn_15_itm_6_rsp_1, NMP_PrepareReadReq_slc_nmp_config_memory_index_1_1_0_itm_7,
      {ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_2_cse , ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_3_cse
      , and_833_nl , and_835_itm , and_836_nl});
  assign ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_not_3_nl = ~ ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_and_1_cse;
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_8_nl
      = MUX_v_2_2_2(2'b00, ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux1h_60_nl,
      ac_math_ac_normalize_40_16_false_AC_TRN_AC_WRAP_expret_not_3_nl);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux1h_59_nl
      = MUX1HOT_v_2_3_2(2'b01, 2'b10, NMP_PrepareWriteReq_slc_nmp_config_memory_index_1_1_0_itm_7,
      {ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_5_cse
      , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_6_cse
      , (~ NMP_RunFSM_switch_lp_conc_itm_7_2)});
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_nand_nl
      = ~((NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z[33:32]==2'b01)
      & NMP_RunFSM_switch_lp_conc_itm_7_2);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_4_nl
      = MUX_v_2_2_2(2'b00, ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_mux1h_59_nl,
      ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_nand_nl);
  assign NMP_PrepareWriteReq_and_nl = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[33:32]==2'b00)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareWriteReq_and_1_nl = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[33:32]==2'b01)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareWriteReq_and_2_nl = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[33:32]==2'b10)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareWriteReq_and_3_nl = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z[33:32]==2'b11)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareWriteReq_NMP_PrepareWriteReq_mux1h_1_nl = MUX1HOT_v_6_4_2(NMP_PrepareWriteReq_asn_1_itm_6_5_0,
      6'b111110, 6'b100110, 6'b110111, {(~ NMP_RunFSM_switch_lp_conc_itm_7_2) , NMP_PrepareWriteReq_and_4_ssc
      , NMP_PrepareWriteReq_and_6_ssc , NMP_PrepareWriteReq_and_7_ssc});
  assign NMP_PrepareWriteReq_not_6_nl = ~ NMP_PrepareWriteReq_and_5_ssc;
  assign NMP_PrepareReadReq_and_2_nl = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[33:32]==2'b00)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareReadReq_and_3_nl = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[33:32]==2'b01)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareReadReq_and_4_nl = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[33:32]==2'b10)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareReadReq_and_5_nl = (NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z[33:32]==2'b11)
      & NMP_RunFSM_switch_lp_conc_itm_7_2;
  assign NMP_PrepareReadReq_NMP_PrepareReadReq_mux1h_1_nl = MUX1HOT_v_6_4_2(NMP_PrepareReadReq_asn_1_itm_6_rsp_1,
      6'b111110, 6'b100110, 6'b110111, {(~ NMP_RunFSM_switch_lp_conc_itm_7_2) , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_7_cse
      , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_5_cse
      , ac_math_ac_pow2_pwl_AC_TRN_33_13_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_output_pwl_and_6_cse});
  assign NMP_PrepareReadReq_not_6_nl = ~ NMP_PrepareReadReq_and_7_ssc;
  assign nmp_config_ConfigRead_nmp_config_ConfigRead_and_7_nl = nmp_config_adpbias_1_sva_mx1_2
      & (~ nmp_config_ConfigRead_unequal_tmp_1);
  assign nmp_config_ConfigRead_not_13_nl = ~ nmp_config_ConfigRead_unequal_tmp_1;
  assign nmp_config_ConfigRead_nmp_config_ConfigRead_and_12_nl = MUX_v_2_2_2(2'b00,
      nmp_config_adpbias_1_sva_mx1_1_0, nmp_config_ConfigRead_not_13_nl);
  assign z_out = MUX_v_8_8_2(8'b00011100, 8'b01001011, 8'b01101100, 8'b10000100,
      8'b10010111, 8'b10100110, 8'b10110011, 8'b10111100, z_out_2[38:36]);
  assign z_out_1 = MUX_v_10_8_2(10'b1111111101, 10'b1100011001, 10'b1001100100, 10'b0111010000,
      10'b0101010100, 10'b0011101011, 10'b0010010001, 10'b0001000100, z_out_2[38:36]);

  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_5_2;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [4:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_5_2;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [4:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    MUX1HOT_v_2_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_5_2;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [4:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    MUX1HOT_v_6_5_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_5_2;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [4:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    MUX1HOT_v_7_5_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input  sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_8_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [2:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_10_8_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [25:0] MUX_v_26_2_2;
    input [25:0] input_0;
    input [25:0] input_1;
    input  sel;
    reg [25:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_26_2_2 = result;
  end
  endfunction


  function automatic [26:0] MUX_v_27_2_2;
    input [26:0] input_0;
    input [26:0] input_1;
    input  sel;
    reg [26:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_27_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [34:0] MUX_v_35_2_2;
    input [34:0] input_0;
    input [34:0] input_1;
    input  sel;
    reg [34:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_35_2_2 = result;
  end
  endfunction


  function automatic [35:0] MUX_v_36_2_2;
    input [35:0] input_0;
    input [35:0] input_1;
    input  sel;
    reg [35:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_36_2_2 = result;
  end
  endfunction


  function automatic [38:0] MUX_v_39_2_2;
    input [38:0] input_0;
    input [38:0] input_1;
    input  sel;
    reg [38:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_39_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_4_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [1:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_3_4_2 = result;
  end
  endfunction


  function automatic [39:0] MUX_v_40_2_2;
    input [39:0] input_0;
    input [39:0] input_1;
    input  sel;
    reg [39:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_40_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_4_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [1:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_5_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_4_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [6:0] input_2;
    input [6:0] input_3;
    input [1:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_7_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_18_1_17;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 17;
    readslicef_18_1_17 = tmp[0:0];
  end
  endfunction


  function automatic [24:0] readslicef_36_25_11;
    input [35:0] vector;
    reg [35:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_36_25_11 = tmp[24:0];
  end
  endfunction


  function automatic [35:0] readslicef_40_36_4;
    input [39:0] vector;
    reg [39:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_40_36_4 = tmp[35:0];
  end
  endfunction


  function automatic [27:0] conv_s2s_27_28 ;
    input [26:0]  vector ;
  begin
    conv_s2s_27_28 = {vector[26], vector};
  end
  endfunction


  function automatic [39:0] conv_s2s_38_40 ;
    input [37:0]  vector ;
  begin
    conv_s2s_38_40 = {{2{vector[37]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2u_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [6:0] conv_s2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2u_6_7 = {vector[5], vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_1_5 ;
    input  vector ;
  begin
    conv_u2s_1_5 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2s_16_18 ;
    input [15:0]  vector ;
  begin
    conv_u2s_16_18 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_1_7 ;
    input  vector ;
  begin
    conv_u2u_1_7 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_9_13 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_13 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction


  function automatic [33:0] conv_u2u_32_34 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_34 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [35:0] conv_u2u_33_36 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_36 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [35:0] conv_u2u_34_36 ;
    input [33:0]  vector ;
  begin
    conv_u2u_34_36 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [36:0] conv_u2u_36_37 ;
    input [35:0]  vector ;
  begin
    conv_u2u_36_37 = {1'b0, vector};
  end
  endfunction


  function automatic [39:0] conv_u2u_39_40 ;
    input [38:0]  vector ;
  begin
    conv_u2u_39_40 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_GBCore
// ------------------------------------------------------------------


module GBModule_GBCore (
  clk, rst, rva_in_large_vld, rva_in_large_rdy, rva_in_large_dat, rva_out_large_vld,
      rva_out_large_rdy, rva_out_large_dat, nmp_large_req_vld, nmp_large_req_rdy,
      nmp_large_req_dat, nmp_large_rsp_vld, nmp_large_rsp_rdy, nmp_large_rsp_dat,
      SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input rva_in_large_vld;
  output rva_in_large_rdy;
  input [168:0] rva_in_large_dat;
  output rva_out_large_vld;
  input rva_out_large_rdy;
  output [127:0] rva_out_large_dat;
  input nmp_large_req_vld;
  output nmp_large_req_rdy;
  input [154:0] nmp_large_req_dat;
  output nmp_large_rsp_vld;
  input nmp_large_rsp_rdy;
  output [127:0] nmp_large_rsp_dat;
  input [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d;
  wire large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a0_a0_a0_a1_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d;
  wire large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a0_a0_a1_a0_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d;
  wire large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a0_a0_a1_a1_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d;
  wire large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a0_a1_a0_a0_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d;
  wire large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a0_a1_a0_a1_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d;
  wire large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a0_a1_a1_a0_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d;
  wire large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a0_a1_a1_a1_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d;
  wire large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a1_a0_a0_a0_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d;
  wire large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a1_a0_a0_a1_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d;
  wire large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a1_a0_a1_a0_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d;
  wire large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a1_a0_a1_a1_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d;
  wire large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a1_a1_a0_a0_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d;
  wire large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a1_a1_a0_a1_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d;
  wire large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a1_a1_a1_a0_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d;
  wire large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d;
  wire [127:0] large_mem_banks_bank_a1_a1_a1_a1_a_rsci_d_d;
  wire [127:0] large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d;
  wire [7:0] GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_a;
  wire [15:0] GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_b;
  wire [11:0] GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_c;
  wire [15:0] GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_z;
  wire large_mem_banks_bank_a0_a0_a0_a0_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsc_q;
  wire large_mem_banks_bank_a0_a0_a0_a0_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsc_radr;
  wire large_mem_banks_bank_a0_a0_a0_a0_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsc_wadr;
  wire large_mem_banks_bank_a0_a0_a0_a1_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a0_a0_a0_a1_a_rsc_q;
  wire large_mem_banks_bank_a0_a0_a0_a1_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a0_a0_a0_a1_a_rsc_radr;
  wire large_mem_banks_bank_a0_a0_a0_a1_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a0_a0_a0_a1_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a0_a0_a0_a1_a_rsc_wadr;
  wire large_mem_banks_bank_a0_a0_a1_a0_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a0_a0_a1_a0_a_rsc_q;
  wire large_mem_banks_bank_a0_a0_a1_a0_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a0_a0_a1_a0_a_rsc_radr;
  wire large_mem_banks_bank_a0_a0_a1_a0_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a0_a0_a1_a0_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a0_a0_a1_a0_a_rsc_wadr;
  wire large_mem_banks_bank_a0_a0_a1_a1_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a0_a0_a1_a1_a_rsc_q;
  wire large_mem_banks_bank_a0_a0_a1_a1_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a0_a0_a1_a1_a_rsc_radr;
  wire large_mem_banks_bank_a0_a0_a1_a1_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a0_a0_a1_a1_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a0_a0_a1_a1_a_rsc_wadr;
  wire large_mem_banks_bank_a0_a1_a0_a0_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a0_a1_a0_a0_a_rsc_q;
  wire large_mem_banks_bank_a0_a1_a0_a0_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a0_a1_a0_a0_a_rsc_radr;
  wire large_mem_banks_bank_a0_a1_a0_a0_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a0_a1_a0_a0_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a0_a1_a0_a0_a_rsc_wadr;
  wire large_mem_banks_bank_a0_a1_a0_a1_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a0_a1_a0_a1_a_rsc_q;
  wire large_mem_banks_bank_a0_a1_a0_a1_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a0_a1_a0_a1_a_rsc_radr;
  wire large_mem_banks_bank_a0_a1_a0_a1_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a0_a1_a0_a1_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a0_a1_a0_a1_a_rsc_wadr;
  wire large_mem_banks_bank_a0_a1_a1_a0_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a0_a1_a1_a0_a_rsc_q;
  wire large_mem_banks_bank_a0_a1_a1_a0_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a0_a1_a1_a0_a_rsc_radr;
  wire large_mem_banks_bank_a0_a1_a1_a0_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a0_a1_a1_a0_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a0_a1_a1_a0_a_rsc_wadr;
  wire large_mem_banks_bank_a0_a1_a1_a1_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a0_a1_a1_a1_a_rsc_q;
  wire large_mem_banks_bank_a0_a1_a1_a1_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a0_a1_a1_a1_a_rsc_radr;
  wire large_mem_banks_bank_a0_a1_a1_a1_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a0_a1_a1_a1_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a0_a1_a1_a1_a_rsc_wadr;
  wire large_mem_banks_bank_a1_a0_a0_a0_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a1_a0_a0_a0_a_rsc_q;
  wire large_mem_banks_bank_a1_a0_a0_a0_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a1_a0_a0_a0_a_rsc_radr;
  wire large_mem_banks_bank_a1_a0_a0_a0_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a1_a0_a0_a0_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a1_a0_a0_a0_a_rsc_wadr;
  wire large_mem_banks_bank_a1_a0_a0_a1_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a1_a0_a0_a1_a_rsc_q;
  wire large_mem_banks_bank_a1_a0_a0_a1_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a1_a0_a0_a1_a_rsc_radr;
  wire large_mem_banks_bank_a1_a0_a0_a1_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a1_a0_a0_a1_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a1_a0_a0_a1_a_rsc_wadr;
  wire large_mem_banks_bank_a1_a0_a1_a0_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a1_a0_a1_a0_a_rsc_q;
  wire large_mem_banks_bank_a1_a0_a1_a0_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a1_a0_a1_a0_a_rsc_radr;
  wire large_mem_banks_bank_a1_a0_a1_a0_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a1_a0_a1_a0_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a1_a0_a1_a0_a_rsc_wadr;
  wire large_mem_banks_bank_a1_a0_a1_a1_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a1_a0_a1_a1_a_rsc_q;
  wire large_mem_banks_bank_a1_a0_a1_a1_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a1_a0_a1_a1_a_rsc_radr;
  wire large_mem_banks_bank_a1_a0_a1_a1_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a1_a0_a1_a1_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a1_a0_a1_a1_a_rsc_wadr;
  wire large_mem_banks_bank_a1_a1_a0_a0_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a1_a1_a0_a0_a_rsc_q;
  wire large_mem_banks_bank_a1_a1_a0_a0_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a1_a1_a0_a0_a_rsc_radr;
  wire large_mem_banks_bank_a1_a1_a0_a0_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a1_a1_a0_a0_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a1_a1_a0_a0_a_rsc_wadr;
  wire large_mem_banks_bank_a1_a1_a0_a1_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a1_a1_a0_a1_a_rsc_q;
  wire large_mem_banks_bank_a1_a1_a0_a1_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a1_a1_a0_a1_a_rsc_radr;
  wire large_mem_banks_bank_a1_a1_a0_a1_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a1_a1_a0_a1_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a1_a1_a0_a1_a_rsc_wadr;
  wire large_mem_banks_bank_a1_a1_a1_a0_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a1_a1_a1_a0_a_rsc_q;
  wire large_mem_banks_bank_a1_a1_a1_a0_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a1_a1_a1_a0_a_rsc_radr;
  wire large_mem_banks_bank_a1_a1_a1_a0_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a1_a1_a1_a0_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a1_a1_a1_a0_a_rsc_wadr;
  wire large_mem_banks_bank_a1_a1_a1_a1_a_rsc_clken;
  wire [127:0] large_mem_banks_bank_a1_a1_a1_a1_a_rsc_q;
  wire large_mem_banks_bank_a1_a1_a1_a1_a_rsc_re;
  wire [11:0] large_mem_banks_bank_a1_a1_a1_a1_a_rsc_radr;
  wire large_mem_banks_bank_a1_a1_a1_a1_a_rsc_we;
  wire [127:0] large_mem_banks_bank_a1_a1_a1_a1_a_rsc_d;
  wire [11:0] large_mem_banks_bank_a1_a1_a1_a1_a_rsc_wadr;
  wire [11:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff;
  wire large_mem_banks_bank_a0_a0_a0_a0_a_rsci_re_d_iff;
  wire [11:0] large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff;
  wire large_mem_banks_bank_a0_a0_a0_a0_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a0_a0_a0_a1_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a0_a0_a0_a1_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a0_a0_a1_a0_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a0_a0_a1_a0_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a0_a0_a1_a1_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a0_a0_a1_a1_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a0_a1_a0_a0_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a0_a1_a0_a0_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a0_a1_a0_a1_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a0_a1_a0_a1_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a0_a1_a1_a0_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a0_a1_a1_a0_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a0_a1_a1_a1_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a0_a1_a1_a1_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a1_a0_a0_a0_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a1_a0_a0_a0_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a1_a0_a0_a1_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a1_a0_a0_a1_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a1_a0_a1_a0_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a1_a0_a1_a0_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a1_a0_a1_a1_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a1_a0_a1_a1_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a1_a1_a0_a0_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a1_a1_a0_a0_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a1_a1_a0_a1_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a1_a1_a0_a1_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a1_a1_a1_a0_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a1_a1_a1_a0_a_rsci_we_d_iff;
  wire large_mem_banks_bank_a1_a1_a1_a1_a_rsci_re_d_iff;
  wire large_mem_banks_bank_a1_a1_a1_a1_a_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_mgc_muladd1 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd12),
  .signd_c(32'sd0),
  .width_cst(32'sd1),
  .signd_cst(32'sd0),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd16),
  .add_axb(32'sd1),
  .add_c(32'sd1),
  .add_d(32'sd1),
  .use_const(32'sd1)) GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp (
      .a(GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_a),
      .b(GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_b),
      .c(GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_c),
      .cst(1'b0),
      .z(GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_z),
      .d(2'b0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a0_a0_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_clken),
      .d(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_d),
      .q(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_q),
      .radr(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_radr),
      .re(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_re),
      .wadr(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_wadr),
      .we(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a0_a0_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_clken),
      .d(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_d),
      .q(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_q),
      .radr(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_radr),
      .re(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_re),
      .wadr(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_wadr),
      .we(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a0_a0_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_clken),
      .d(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_d),
      .q(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_q),
      .radr(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_radr),
      .re(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_re),
      .wadr(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_wadr),
      .we(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a0_a0_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_clken),
      .d(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_d),
      .q(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_q),
      .radr(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_radr),
      .re(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_re),
      .wadr(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_wadr),
      .we(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a0_a1_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_clken),
      .d(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_d),
      .q(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_q),
      .radr(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_radr),
      .re(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_re),
      .wadr(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_wadr),
      .we(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a0_a1_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_clken),
      .d(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_d),
      .q(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_q),
      .radr(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_radr),
      .re(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_re),
      .wadr(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_wadr),
      .we(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a0_a1_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_clken),
      .d(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_d),
      .q(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_q),
      .radr(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_radr),
      .re(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_re),
      .wadr(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_wadr),
      .we(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a0_a1_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_clken),
      .d(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_d),
      .q(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_q),
      .radr(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_radr),
      .re(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_re),
      .wadr(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_wadr),
      .we(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a1_a0_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_clken),
      .d(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_d),
      .q(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_q),
      .radr(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_radr),
      .re(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_re),
      .wadr(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_wadr),
      .we(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a1_a0_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_clken),
      .d(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_d),
      .q(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_q),
      .radr(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_radr),
      .re(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_re),
      .wadr(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_wadr),
      .we(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a1_a0_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_clken),
      .d(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_d),
      .q(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_q),
      .radr(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_radr),
      .re(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_re),
      .wadr(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_wadr),
      .we(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a1_a0_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_clken),
      .d(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_d),
      .q(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_q),
      .radr(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_radr),
      .re(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_re),
      .wadr(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_wadr),
      .we(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a1_a1_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_clken),
      .d(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_d),
      .q(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_q),
      .radr(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_radr),
      .re(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_re),
      .wadr(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_wadr),
      .we(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a1_a1_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_clken),
      .d(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_d),
      .q(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_q),
      .radr(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_radr),
      .re(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_re),
      .wadr(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_wadr),
      .we(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a1_a1_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_clken),
      .d(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_d),
      .q(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_q),
      .radr(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_radr),
      .re(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_re),
      .wadr(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_wadr),
      .we(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) large_mem_banks_bank_a1_a1_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_clken),
      .d(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_d),
      .q(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_q),
      .radr(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_radr),
      .re(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_re),
      .wadr(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_wadr),
      .we(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_we)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_62_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a0_a0_a0_a0_a_rsci (
      .clken(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_clken),
      .q(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_q),
      .re(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_re),
      .radr(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_radr),
      .we(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_we),
      .d(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_d),
      .wadr(large_mem_banks_bank_a0_a0_a0_a0_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_63_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a0_a0_a0_a1_a_rsci (
      .clken(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_clken),
      .q(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_q),
      .re(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_re),
      .radr(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_radr),
      .we(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_we),
      .d(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_d),
      .wadr(large_mem_banks_bank_a0_a0_a0_a1_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_64_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a0_a0_a1_a0_a_rsci (
      .clken(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_clken),
      .q(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_q),
      .re(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_re),
      .radr(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_radr),
      .we(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_we),
      .d(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_d),
      .wadr(large_mem_banks_bank_a0_a0_a1_a0_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_65_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a0_a0_a1_a1_a_rsci (
      .clken(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_clken),
      .q(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_q),
      .re(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_re),
      .radr(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_radr),
      .we(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_we),
      .d(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_d),
      .wadr(large_mem_banks_bank_a0_a0_a1_a1_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_66_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a0_a1_a0_a0_a_rsci (
      .clken(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_clken),
      .q(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_q),
      .re(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_re),
      .radr(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_radr),
      .we(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_we),
      .d(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_d),
      .wadr(large_mem_banks_bank_a0_a1_a0_a0_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_67_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a0_a1_a0_a1_a_rsci (
      .clken(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_clken),
      .q(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_q),
      .re(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_re),
      .radr(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_radr),
      .we(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_we),
      .d(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_d),
      .wadr(large_mem_banks_bank_a0_a1_a0_a1_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_68_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a0_a1_a1_a0_a_rsci (
      .clken(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_clken),
      .q(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_q),
      .re(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_re),
      .radr(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_radr),
      .we(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_we),
      .d(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_d),
      .wadr(large_mem_banks_bank_a0_a1_a1_a0_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_69_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a0_a1_a1_a1_a_rsci (
      .clken(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_clken),
      .q(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_q),
      .re(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_re),
      .radr(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_radr),
      .we(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_we),
      .d(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_d),
      .wadr(large_mem_banks_bank_a0_a1_a1_a1_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_70_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a1_a0_a0_a0_a_rsci (
      .clken(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_clken),
      .q(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_q),
      .re(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_re),
      .radr(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_radr),
      .we(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_we),
      .d(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_d),
      .wadr(large_mem_banks_bank_a1_a0_a0_a0_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_71_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a1_a0_a0_a1_a_rsci (
      .clken(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_clken),
      .q(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_q),
      .re(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_re),
      .radr(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_radr),
      .we(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_we),
      .d(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_d),
      .wadr(large_mem_banks_bank_a1_a0_a0_a1_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_72_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a1_a0_a1_a0_a_rsci (
      .clken(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_clken),
      .q(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_q),
      .re(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_re),
      .radr(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_radr),
      .we(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_we),
      .d(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_d),
      .wadr(large_mem_banks_bank_a1_a0_a1_a0_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_73_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a1_a0_a1_a1_a_rsci (
      .clken(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_clken),
      .q(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_q),
      .re(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_re),
      .radr(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_radr),
      .we(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_we),
      .d(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_d),
      .wadr(large_mem_banks_bank_a1_a0_a1_a1_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_74_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a1_a1_a0_a0_a_rsci (
      .clken(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_clken),
      .q(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_q),
      .re(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_re),
      .radr(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_radr),
      .we(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_we),
      .d(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_d),
      .wadr(large_mem_banks_bank_a1_a1_a0_a0_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_75_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a1_a1_a0_a1_a_rsci (
      .clken(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_clken),
      .q(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_q),
      .re(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_re),
      .radr(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_radr),
      .we(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_we),
      .d(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_d),
      .wadr(large_mem_banks_bank_a1_a1_a0_a1_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_76_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a1_a1_a1_a0_a_rsci (
      .clken(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_clken),
      .q(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_q),
      .re(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_re),
      .radr(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_radr),
      .we(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_we),
      .d(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_d),
      .wadr(large_mem_banks_bank_a1_a1_a1_a0_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_re_d_iff)
    );
  GBModule_GBCore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_77_12_128_4096_1_4096_128_1_gen
      large_mem_banks_bank_a1_a1_a1_a1_a_rsci (
      .clken(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_clken),
      .q(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_q),
      .re(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_re),
      .radr(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_radr),
      .we(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_we),
      .d(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_d),
      .wadr(large_mem_banks_bank_a1_a1_a1_a1_a_rsc_wadr),
      .clken_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d),
      .d_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_d_d),
      .q_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d),
      .radr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .re_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_re_d_iff),
      .wadr_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_re_d_iff)
    );
  GBModule_GBCore_GBCoreRun GBCore_GBCoreRun_inst (
      .clk(clk),
      .rst(rst),
      .rva_in_large_vld(rva_in_large_vld),
      .rva_in_large_rdy(rva_in_large_rdy),
      .rva_in_large_dat(rva_in_large_dat),
      .rva_out_large_vld(rva_out_large_vld),
      .rva_out_large_rdy(rva_out_large_rdy),
      .rva_out_large_dat(rva_out_large_dat),
      .nmp_large_req_vld(nmp_large_req_vld),
      .nmp_large_req_rdy(nmp_large_req_rdy),
      .nmp_large_req_dat(nmp_large_req_dat),
      .nmp_large_rsp_vld(nmp_large_rsp_vld),
      .nmp_large_rsp_rdy(nmp_large_rsp_rdy),
      .nmp_large_rsp_dat(nmp_large_rsp_dat),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG),
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_d_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_d_d),
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_q_d),
      .large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a0_a0_a1_a_rsci_d_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_d_d),
      .large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_q_d),
      .large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a0_a1_a0_a_rsci_d_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_d_d),
      .large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_q_d),
      .large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a0_a1_a1_a_rsci_d_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_d_d),
      .large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_q_d),
      .large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a1_a0_a0_a_rsci_d_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_d_d),
      .large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_q_d),
      .large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a1_a0_a1_a_rsci_d_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_d_d),
      .large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_q_d),
      .large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a1_a1_a0_a_rsci_d_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_d_d),
      .large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_q_d),
      .large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a0_a1_a1_a1_a_rsci_d_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_d_d),
      .large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_q_d),
      .large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a0_a0_a0_a_rsci_d_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_d_d),
      .large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_q_d),
      .large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a0_a0_a1_a_rsci_d_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_d_d),
      .large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_q_d),
      .large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a0_a1_a0_a_rsci_d_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_d_d),
      .large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_q_d),
      .large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a0_a1_a1_a_rsci_d_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_d_d),
      .large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_q_d),
      .large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a1_a0_a0_a_rsci_d_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_d_d),
      .large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_q_d),
      .large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a1_a0_a1_a_rsci_d_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_d_d),
      .large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_q_d),
      .large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a1_a1_a0_a_rsci_d_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_d_d),
      .large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_q_d),
      .large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_clken_d),
      .large_mem_banks_bank_a1_a1_a1_a1_a_rsci_d_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_d_d),
      .large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_q_d),
      .GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_a(GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_a),
      .GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_b(GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_b),
      .GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_c(GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_c),
      .GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_z(GBCore_SetLargeBuffer_1U_base_addr_acc_4_cmp_z),
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_pff(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_radr_d_iff),
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_re_d_pff(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_re_d_iff),
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_pff(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_wadr_d_iff),
      .large_mem_banks_bank_a0_a0_a0_a0_a_rsci_we_d_pff(large_mem_banks_bank_a0_a0_a0_a0_a_rsci_we_d_iff),
      .large_mem_banks_bank_a0_a0_a0_a1_a_rsci_re_d_pff(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_re_d_iff),
      .large_mem_banks_bank_a0_a0_a0_a1_a_rsci_we_d_pff(large_mem_banks_bank_a0_a0_a0_a1_a_rsci_we_d_iff),
      .large_mem_banks_bank_a0_a0_a1_a0_a_rsci_re_d_pff(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_re_d_iff),
      .large_mem_banks_bank_a0_a0_a1_a0_a_rsci_we_d_pff(large_mem_banks_bank_a0_a0_a1_a0_a_rsci_we_d_iff),
      .large_mem_banks_bank_a0_a0_a1_a1_a_rsci_re_d_pff(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_re_d_iff),
      .large_mem_banks_bank_a0_a0_a1_a1_a_rsci_we_d_pff(large_mem_banks_bank_a0_a0_a1_a1_a_rsci_we_d_iff),
      .large_mem_banks_bank_a0_a1_a0_a0_a_rsci_re_d_pff(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_re_d_iff),
      .large_mem_banks_bank_a0_a1_a0_a0_a_rsci_we_d_pff(large_mem_banks_bank_a0_a1_a0_a0_a_rsci_we_d_iff),
      .large_mem_banks_bank_a0_a1_a0_a1_a_rsci_re_d_pff(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_re_d_iff),
      .large_mem_banks_bank_a0_a1_a0_a1_a_rsci_we_d_pff(large_mem_banks_bank_a0_a1_a0_a1_a_rsci_we_d_iff),
      .large_mem_banks_bank_a0_a1_a1_a0_a_rsci_re_d_pff(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_re_d_iff),
      .large_mem_banks_bank_a0_a1_a1_a0_a_rsci_we_d_pff(large_mem_banks_bank_a0_a1_a1_a0_a_rsci_we_d_iff),
      .large_mem_banks_bank_a0_a1_a1_a1_a_rsci_re_d_pff(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_re_d_iff),
      .large_mem_banks_bank_a0_a1_a1_a1_a_rsci_we_d_pff(large_mem_banks_bank_a0_a1_a1_a1_a_rsci_we_d_iff),
      .large_mem_banks_bank_a1_a0_a0_a0_a_rsci_re_d_pff(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_re_d_iff),
      .large_mem_banks_bank_a1_a0_a0_a0_a_rsci_we_d_pff(large_mem_banks_bank_a1_a0_a0_a0_a_rsci_we_d_iff),
      .large_mem_banks_bank_a1_a0_a0_a1_a_rsci_re_d_pff(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_re_d_iff),
      .large_mem_banks_bank_a1_a0_a0_a1_a_rsci_we_d_pff(large_mem_banks_bank_a1_a0_a0_a1_a_rsci_we_d_iff),
      .large_mem_banks_bank_a1_a0_a1_a0_a_rsci_re_d_pff(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_re_d_iff),
      .large_mem_banks_bank_a1_a0_a1_a0_a_rsci_we_d_pff(large_mem_banks_bank_a1_a0_a1_a0_a_rsci_we_d_iff),
      .large_mem_banks_bank_a1_a0_a1_a1_a_rsci_re_d_pff(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_re_d_iff),
      .large_mem_banks_bank_a1_a0_a1_a1_a_rsci_we_d_pff(large_mem_banks_bank_a1_a0_a1_a1_a_rsci_we_d_iff),
      .large_mem_banks_bank_a1_a1_a0_a0_a_rsci_re_d_pff(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_re_d_iff),
      .large_mem_banks_bank_a1_a1_a0_a0_a_rsci_we_d_pff(large_mem_banks_bank_a1_a1_a0_a0_a_rsci_we_d_iff),
      .large_mem_banks_bank_a1_a1_a0_a1_a_rsci_re_d_pff(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_re_d_iff),
      .large_mem_banks_bank_a1_a1_a0_a1_a_rsci_we_d_pff(large_mem_banks_bank_a1_a1_a0_a1_a_rsci_we_d_iff),
      .large_mem_banks_bank_a1_a1_a1_a0_a_rsci_re_d_pff(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_re_d_iff),
      .large_mem_banks_bank_a1_a1_a1_a0_a_rsci_we_d_pff(large_mem_banks_bank_a1_a1_a1_a0_a_rsci_we_d_iff),
      .large_mem_banks_bank_a1_a1_a1_a1_a_rsci_re_d_pff(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_re_d_iff),
      .large_mem_banks_bank_a1_a1_a1_a1_a_rsci_we_d_pff(large_mem_banks_bank_a1_a1_a1_a1_a_rsci_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule_NMP
// ------------------------------------------------------------------


module GBModule_NMP (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      start_vld, start_rdy, start_dat, done_vld, done_rdy, done_dat, large_req_vld,
      large_req_rdy, large_req_dat, large_rsp_vld, large_rsp_rdy, large_rsp_dat
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  input start_vld;
  output start_rdy;
  input start_dat;
  output done_vld;
  input done_rdy;
  output done_dat;
  output large_req_vld;
  input large_req_rdy;
  output [154:0] large_req_dat;
  input large_rsp_vld;
  output large_rsp_rdy;
  input [127:0] large_rsp_dat;


  // Interconnect Declarations
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_a;
  wire NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_z;
  wire [31:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_a;
  wire [55:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_b;
  wire NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z;
  wire [27:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_b;
  wire [42:0] NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_a;
  wire NMP_ComputeRMSNormalize_for_1_mul_cmp_en;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_1_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_1_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_2_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_2_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_3_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_3_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_4_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_4_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_5_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_5_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_6_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_6_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_7_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_7_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_8_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_8_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_9_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_9_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_10_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_10_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_11_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_11_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_12_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_12_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_13_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_13_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_14_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_14_z;
  wire [26:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_15_a;
  wire [55:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_15_z;
  wire NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_z;
  wire [53:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_z;
  wire [39:0] NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff;
  wire [39:0] NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_a_iff;
  wire [26:0] NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_a_iff;


  // Interconnect Declarations for Component Instantiations 
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15 (
      .a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_a),
      .b(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_b(32'sd28),
  .signd_b(32'sd1),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15
      (
      .a(15'b101110001010101),
      .b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_b),
      .clk(clk),
      .en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_1 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_1_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_1_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_2 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_2_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_2_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_3 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_3_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_3_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_4 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_4_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_4_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_5 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_5_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_5_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_6 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_6_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_6_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_7 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_7_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_7_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_8 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_8_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_8_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_9 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_9_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_9_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_10 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_10_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_10_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_11 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_11_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_11_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_12 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_12_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_12_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_13 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_13_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_13_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_14 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_14_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_14_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd40),
  .signd_b(32'sd1),
  .width_z(32'sd56),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) NMP_ComputeRMSNormalize_for_1_mul_cmp_15 (
      .a(NMP_ComputeRMSNormalize_for_1_mul_cmp_15_a),
      .b(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .clk(clk),
      .en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSNormalize_for_1_mul_cmp_15_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1 (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2 (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3 (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4 (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5 (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6 (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7 (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8 (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9 (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10
      (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11
      (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12
      (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13
      (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14
      (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_z)
    );
  GBModule_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15
      (
      .a(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_a_iff),
      .b(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_a_iff),
      .clk(clk),
      .en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_z)
    );
  GBModule_NMP_NMPRun NMP_NMPRun_inst (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .done_vld(done_vld),
      .done_rdy(done_rdy),
      .done_dat(done_dat),
      .large_req_vld(large_req_vld),
      .large_req_rdy(large_req_rdy),
      .large_req_dat(large_req_dat),
      .large_rsp_vld(large_rsp_vld),
      .large_rsp_rdy(large_rsp_rdy),
      .large_rsp_dat(large_rsp_dat),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_en),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_1_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_2_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_3_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_4_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_5_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_6_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_7_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_8_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_9_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_10_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_11_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_12_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_13_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_14_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_a(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_a),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_z(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_15_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_en),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_1_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_2_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_3_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_4_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_5_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_6_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_7_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_8_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_9_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_10_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_11_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_12_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_13_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_14_z),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_b(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_b),
      .NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z(NMP_ComputeSoftmaxExp_for_1_ac_math_ac_exp_pwl_11_AC_TRN_32_12_true_AC_TRN_AC_WRAP_32_12_AC_TRN_AC_WRAP_mul_cmp_15_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_en(NMP_ComputeRMSNormalize_for_1_mul_cmp_en),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_1_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_1_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_1_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_1_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_2_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_2_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_2_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_2_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_3_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_3_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_3_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_3_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_4_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_4_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_4_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_4_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_5_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_5_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_5_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_5_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_6_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_6_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_6_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_6_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_7_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_7_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_7_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_7_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_8_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_8_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_8_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_8_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_9_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_9_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_9_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_9_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_10_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_10_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_10_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_10_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_11_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_11_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_11_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_11_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_12_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_12_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_12_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_12_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_13_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_13_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_13_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_13_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_14_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_14_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_14_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_14_z),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_15_a(NMP_ComputeRMSNormalize_for_1_mul_cmp_15_a),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_15_z(NMP_ComputeRMSNormalize_for_1_mul_cmp_15_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_en),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_z),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_z(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_z),
      .NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_pff(NMP_ComputeSoftmaxNormalize_for_1_mul_cmp_b_iff),
      .NMP_ComputeRMSNormalize_for_1_mul_cmp_b_pff(NMP_ComputeRMSNormalize_for_1_mul_cmp_b_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_1_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_2_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_3_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_4_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_5_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_6_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_7_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_8_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_9_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_10_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_11_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_12_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_13_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_14_a_iff),
      .NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_a_pff(NMP_ComputeRMSSumSq_for_1_NMP_ComputeRMSSumSq_for_mul_cmp_15_a_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    GBModule
// ------------------------------------------------------------------


module GBModule (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      start_vld, start_rdy, start_dat, done_vld, done_rdy, done_dat
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  input start_vld;
  output start_rdy;
  input start_dat;
  output done_vld;
  input done_rdy;
  output done_dat;


  // Interconnect Declarations
  wire gbcore_rva_in_vld;
  wire gbcore_rva_in_rdy;
  wire [168:0] gbcore_rva_in_dat;
  wire gbcore_rva_out_vld;
  wire gbcore_rva_out_rdy;
  wire [127:0] gbcore_rva_out_dat;
  wire nmp_rva_in_vld;
  wire nmp_rva_in_rdy;
  wire [168:0] nmp_rva_in_dat;
  wire nmp_rva_out_vld;
  wire nmp_rva_out_rdy;
  wire [127:0] nmp_rva_out_dat;
  wire nmp_large_req_vld;
  wire nmp_large_req_rdy;
  wire [154:0] nmp_large_req_dat;
  wire nmp_large_rsp_vld;
  wire nmp_large_rsp_rdy;
  wire [127:0] nmp_large_rsp_dat;
  wire [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations for Component Instantiations 
  GBModule_GBCore gbcore_inst (
      .clk(clk),
      .rst(rst),
      .rva_in_large_vld(gbcore_rva_in_vld),
      .rva_in_large_rdy(gbcore_rva_in_rdy),
      .rva_in_large_dat(gbcore_rva_in_dat),
      .rva_out_large_vld(gbcore_rva_out_vld),
      .rva_out_large_rdy(gbcore_rva_out_rdy),
      .rva_out_large_dat(gbcore_rva_out_dat),
      .nmp_large_req_vld(nmp_large_req_vld),
      .nmp_large_req_rdy(nmp_large_req_rdy),
      .nmp_large_req_dat(nmp_large_req_dat),
      .nmp_large_rsp_vld(nmp_large_rsp_vld),
      .nmp_large_rsp_rdy(nmp_large_rsp_rdy),
      .nmp_large_rsp_dat(nmp_large_rsp_dat),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG)
    );
  GBModule_NMP nmp_inst (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(nmp_rva_in_vld),
      .rva_in_rdy(nmp_rva_in_rdy),
      .rva_in_dat(nmp_rva_in_dat),
      .rva_out_vld(nmp_rva_out_vld),
      .rva_out_rdy(nmp_rva_out_rdy),
      .rva_out_dat(nmp_rva_out_dat),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .done_vld(done_vld),
      .done_rdy(done_rdy),
      .done_dat(done_dat),
      .large_req_vld(nmp_large_req_vld),
      .large_req_rdy(nmp_large_req_rdy),
      .large_req_dat(nmp_large_req_dat),
      .large_rsp_vld(nmp_large_rsp_vld),
      .large_rsp_rdy(nmp_large_rsp_rdy),
      .large_rsp_dat(nmp_large_rsp_dat)
    );
  GBModule_GBModule_RVAInRun GBModule_RVAInRun_inst (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .gbcore_rva_in_vld(gbcore_rva_in_vld),
      .gbcore_rva_in_rdy(gbcore_rva_in_rdy),
      .gbcore_rva_in_dat(gbcore_rva_in_dat),
      .nmp_rva_in_vld(nmp_rva_in_vld),
      .nmp_rva_in_rdy(nmp_rva_in_rdy),
      .nmp_rva_in_dat(nmp_rva_in_dat),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG)
    );
  GBModule_GBModule_RVAOutRun GBModule_RVAOutRun_inst (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .gbcore_rva_out_vld(gbcore_rva_out_vld),
      .gbcore_rva_out_rdy(gbcore_rva_out_rdy),
      .gbcore_rva_out_dat(gbcore_rva_out_dat),
      .nmp_rva_out_vld(nmp_rva_out_vld),
      .nmp_rva_out_rdy(nmp_rva_out_rdy),
      .nmp_rva_out_dat(nmp_rva_out_dat)
    );
endmodule



